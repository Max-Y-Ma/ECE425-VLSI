* SPICE NETLIST
***************************************

.SUBCKT M1_POLY_CDNS_712253429492
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NTAP_CDNS_712253429491
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PTAP_CDNS_712253429490
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=3 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172
** N=1092 EP=172 IP=2241 FDC=2700
M0 173 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=134870 $D=1
M1 174 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=139500 $D=1
M2 175 1 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=144130 $D=1
M3 176 173 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=134870 $D=1
M4 177 174 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=139500 $D=1
M5 178 175 4 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=144130 $D=1
M6 8 1 176 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=134870 $D=1
M7 9 1 177 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=139500 $D=1
M8 140 1 178 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=144130 $D=1
M9 179 173 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=134870 $D=1
M10 180 174 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=139500 $D=1
M11 181 175 4 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=144130 $D=1
M12 2 1 179 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=134870 $D=1
M13 3 1 180 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=139500 $D=1
M14 4 1 181 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=144130 $D=1
M15 182 173 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=134870 $D=1
M16 183 174 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=139500 $D=1
M17 184 175 4 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=144130 $D=1
M18 2 1 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=134870 $D=1
M19 3 1 183 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=139500 $D=1
M20 4 1 184 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=144130 $D=1
M21 188 185 182 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=134870 $D=1
M22 189 186 183 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=139500 $D=1
M23 190 187 184 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=144130 $D=1
M24 185 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=134870 $D=1
M25 186 5 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=139500 $D=1
M26 187 5 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=144130 $D=1
M27 191 185 179 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=134870 $D=1
M28 192 186 180 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=139500 $D=1
M29 193 187 181 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=144130 $D=1
M30 176 5 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=134870 $D=1
M31 177 5 192 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=139500 $D=1
M32 178 5 193 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=144130 $D=1
M33 194 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=134870 $D=1
M34 195 6 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=139500 $D=1
M35 196 6 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=144130 $D=1
M36 197 194 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=134870 $D=1
M37 198 195 192 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=139500 $D=1
M38 199 196 193 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=144130 $D=1
M39 188 6 197 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=134870 $D=1
M40 189 6 198 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=139500 $D=1
M41 190 6 199 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=144130 $D=1
M42 200 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=134870 $D=1
M43 201 7 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=139500 $D=1
M44 202 7 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=144130 $D=1
M45 203 200 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=134870 $D=1
M46 204 201 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=139500 $D=1
M47 205 202 10 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=144130 $D=1
M48 11 7 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=134870 $D=1
M49 12 7 204 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=139500 $D=1
M50 13 7 205 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=144130 $D=1
M51 206 200 14 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=134870 $D=1
M52 207 201 15 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=139500 $D=1
M53 208 202 16 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=144130 $D=1
M54 209 7 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=134870 $D=1
M55 210 7 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=139500 $D=1
M56 211 7 208 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=144130 $D=1
M57 215 200 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=134870 $D=1
M58 216 201 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=139500 $D=1
M59 217 202 214 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=144130 $D=1
M60 197 7 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=134870 $D=1
M61 198 7 216 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=139500 $D=1
M62 199 7 217 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=144130 $D=1
M63 221 218 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=134870 $D=1
M64 222 219 216 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=139500 $D=1
M65 223 220 217 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=144130 $D=1
M66 218 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=134870 $D=1
M67 219 17 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=139500 $D=1
M68 220 17 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=144130 $D=1
M69 224 218 206 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=134870 $D=1
M70 225 219 207 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=139500 $D=1
M71 226 220 208 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=144130 $D=1
M72 203 17 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=134870 $D=1
M73 204 17 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=139500 $D=1
M74 205 17 226 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=144130 $D=1
M75 227 18 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=134870 $D=1
M76 228 18 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=139500 $D=1
M77 229 18 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=144130 $D=1
M78 230 227 224 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=134870 $D=1
M79 231 228 225 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=139500 $D=1
M80 232 229 226 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=144130 $D=1
M81 221 18 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=134870 $D=1
M82 222 18 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=139500 $D=1
M83 223 18 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=144130 $D=1
M84 8 19 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=134870 $D=1
M85 9 19 234 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=139500 $D=1
M86 140 19 235 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=144130 $D=1
M87 236 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=134870 $D=1
M88 237 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=139500 $D=1
M89 238 20 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=144130 $D=1
M90 239 19 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=134870 $D=1
M91 240 19 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=139500 $D=1
M92 241 19 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=144130 $D=1
M93 8 239 940 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=134870 $D=1
M94 9 240 941 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=139500 $D=1
M95 140 241 942 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=144130 $D=1
M96 242 940 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=134870 $D=1
M97 243 941 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=139500 $D=1
M98 244 942 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=144130 $D=1
M99 239 233 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=134870 $D=1
M100 240 234 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=139500 $D=1
M101 241 235 244 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=144130 $D=1
M102 242 20 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=134870 $D=1
M103 243 20 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=139500 $D=1
M104 244 20 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=144130 $D=1
M105 251 21 242 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=134870 $D=1
M106 252 21 243 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=139500 $D=1
M107 253 21 244 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=144130 $D=1
M108 248 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=134870 $D=1
M109 249 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=139500 $D=1
M110 250 21 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=144130 $D=1
M111 8 22 254 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=134870 $D=1
M112 9 22 255 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=139500 $D=1
M113 140 22 256 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=144130 $D=1
M114 257 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=134870 $D=1
M115 258 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=139500 $D=1
M116 259 23 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=144130 $D=1
M117 260 22 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=134870 $D=1
M118 261 22 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=139500 $D=1
M119 262 22 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=144130 $D=1
M120 8 260 943 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=134870 $D=1
M121 9 261 944 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=139500 $D=1
M122 140 262 945 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=144130 $D=1
M123 263 943 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=134870 $D=1
M124 264 944 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=139500 $D=1
M125 265 945 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=144130 $D=1
M126 260 254 263 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=134870 $D=1
M127 261 255 264 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=139500 $D=1
M128 262 256 265 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=144130 $D=1
M129 263 23 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=134870 $D=1
M130 264 23 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=139500 $D=1
M131 265 23 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=144130 $D=1
M132 251 24 263 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=134870 $D=1
M133 252 24 264 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=139500 $D=1
M134 253 24 265 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=144130 $D=1
M135 266 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=134870 $D=1
M136 267 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=139500 $D=1
M137 268 24 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=144130 $D=1
M138 8 25 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=134870 $D=1
M139 9 25 270 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=139500 $D=1
M140 140 25 271 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=144130 $D=1
M141 272 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=134870 $D=1
M142 273 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=139500 $D=1
M143 274 26 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=144130 $D=1
M144 275 25 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=134870 $D=1
M145 276 25 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=139500 $D=1
M146 277 25 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=144130 $D=1
M147 8 275 946 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=134870 $D=1
M148 9 276 947 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=139500 $D=1
M149 140 277 948 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=144130 $D=1
M150 278 946 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=134870 $D=1
M151 279 947 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=139500 $D=1
M152 280 948 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=144130 $D=1
M153 275 269 278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=134870 $D=1
M154 276 270 279 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=139500 $D=1
M155 277 271 280 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=144130 $D=1
M156 278 26 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=134870 $D=1
M157 279 26 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=139500 $D=1
M158 280 26 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=144130 $D=1
M159 251 27 278 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=134870 $D=1
M160 252 27 279 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=139500 $D=1
M161 253 27 280 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=144130 $D=1
M162 281 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=134870 $D=1
M163 282 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=139500 $D=1
M164 283 27 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=144130 $D=1
M165 8 28 284 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=134870 $D=1
M166 9 28 285 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=139500 $D=1
M167 140 28 286 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=144130 $D=1
M168 287 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=134870 $D=1
M169 288 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=139500 $D=1
M170 289 29 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=144130 $D=1
M171 290 28 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=134870 $D=1
M172 291 28 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=139500 $D=1
M173 292 28 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=144130 $D=1
M174 8 290 949 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=134870 $D=1
M175 9 291 950 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=139500 $D=1
M176 140 292 951 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=144130 $D=1
M177 293 949 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=134870 $D=1
M178 294 950 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=139500 $D=1
M179 295 951 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=144130 $D=1
M180 290 284 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=134870 $D=1
M181 291 285 294 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=139500 $D=1
M182 292 286 295 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=144130 $D=1
M183 293 29 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=134870 $D=1
M184 294 29 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=139500 $D=1
M185 295 29 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=144130 $D=1
M186 251 30 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=134870 $D=1
M187 252 30 294 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=139500 $D=1
M188 253 30 295 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=144130 $D=1
M189 296 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=134870 $D=1
M190 297 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=139500 $D=1
M191 298 30 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=144130 $D=1
M192 8 31 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=134870 $D=1
M193 9 31 300 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=139500 $D=1
M194 140 31 301 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=144130 $D=1
M195 302 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=134870 $D=1
M196 303 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=139500 $D=1
M197 304 32 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=144130 $D=1
M198 305 31 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=134870 $D=1
M199 306 31 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=139500 $D=1
M200 307 31 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=144130 $D=1
M201 8 305 952 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=134870 $D=1
M202 9 306 953 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=139500 $D=1
M203 140 307 954 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=144130 $D=1
M204 308 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=134870 $D=1
M205 309 953 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=139500 $D=1
M206 310 954 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=144130 $D=1
M207 305 299 308 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=134870 $D=1
M208 306 300 309 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=139500 $D=1
M209 307 301 310 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=144130 $D=1
M210 308 32 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=134870 $D=1
M211 309 32 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=139500 $D=1
M212 310 32 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=144130 $D=1
M213 251 33 308 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=134870 $D=1
M214 252 33 309 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=139500 $D=1
M215 253 33 310 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=144130 $D=1
M216 311 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=134870 $D=1
M217 312 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=139500 $D=1
M218 313 33 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=144130 $D=1
M219 8 34 314 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=134870 $D=1
M220 9 34 315 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=139500 $D=1
M221 140 34 316 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=144130 $D=1
M222 317 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=134870 $D=1
M223 318 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=139500 $D=1
M224 319 35 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=144130 $D=1
M225 320 34 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=134870 $D=1
M226 321 34 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=139500 $D=1
M227 322 34 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=144130 $D=1
M228 8 320 955 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=134870 $D=1
M229 9 321 956 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=139500 $D=1
M230 140 322 957 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=144130 $D=1
M231 323 955 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=134870 $D=1
M232 324 956 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=139500 $D=1
M233 325 957 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=144130 $D=1
M234 320 314 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=134870 $D=1
M235 321 315 324 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=139500 $D=1
M236 322 316 325 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=144130 $D=1
M237 323 35 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=134870 $D=1
M238 324 35 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=139500 $D=1
M239 325 35 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=144130 $D=1
M240 251 36 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=134870 $D=1
M241 252 36 324 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=139500 $D=1
M242 253 36 325 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=144130 $D=1
M243 326 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=134870 $D=1
M244 327 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=139500 $D=1
M245 328 36 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=144130 $D=1
M246 8 37 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=134870 $D=1
M247 9 37 330 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=139500 $D=1
M248 140 37 331 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=144130 $D=1
M249 332 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=134870 $D=1
M250 333 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=139500 $D=1
M251 334 38 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=144130 $D=1
M252 335 37 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=134870 $D=1
M253 336 37 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=139500 $D=1
M254 337 37 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=144130 $D=1
M255 8 335 958 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=134870 $D=1
M256 9 336 959 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=139500 $D=1
M257 140 337 960 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=144130 $D=1
M258 338 958 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=134870 $D=1
M259 339 959 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=139500 $D=1
M260 340 960 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=144130 $D=1
M261 335 329 338 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=134870 $D=1
M262 336 330 339 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=139500 $D=1
M263 337 331 340 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=144130 $D=1
M264 338 38 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=134870 $D=1
M265 339 38 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=139500 $D=1
M266 340 38 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=144130 $D=1
M267 251 39 338 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=134870 $D=1
M268 252 39 339 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=139500 $D=1
M269 253 39 340 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=144130 $D=1
M270 341 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=134870 $D=1
M271 342 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=139500 $D=1
M272 343 39 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=144130 $D=1
M273 8 40 344 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=134870 $D=1
M274 9 40 345 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=139500 $D=1
M275 140 40 346 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=144130 $D=1
M276 347 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=134870 $D=1
M277 348 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=139500 $D=1
M278 349 41 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=144130 $D=1
M279 350 40 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=134870 $D=1
M280 351 40 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=139500 $D=1
M281 352 40 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=144130 $D=1
M282 8 350 961 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=134870 $D=1
M283 9 351 962 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=139500 $D=1
M284 140 352 963 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=144130 $D=1
M285 353 961 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=134870 $D=1
M286 354 962 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=139500 $D=1
M287 355 963 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=144130 $D=1
M288 350 344 353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=134870 $D=1
M289 351 345 354 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=139500 $D=1
M290 352 346 355 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=144130 $D=1
M291 353 41 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=134870 $D=1
M292 354 41 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=139500 $D=1
M293 355 41 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=144130 $D=1
M294 251 42 353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=134870 $D=1
M295 252 42 354 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=139500 $D=1
M296 253 42 355 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=144130 $D=1
M297 356 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=134870 $D=1
M298 357 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=139500 $D=1
M299 358 42 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=144130 $D=1
M300 8 43 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=134870 $D=1
M301 9 43 360 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=139500 $D=1
M302 140 43 361 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=144130 $D=1
M303 362 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=134870 $D=1
M304 363 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=139500 $D=1
M305 364 44 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=144130 $D=1
M306 365 43 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=134870 $D=1
M307 366 43 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=139500 $D=1
M308 367 43 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=144130 $D=1
M309 8 365 964 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=134870 $D=1
M310 9 366 965 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=139500 $D=1
M311 140 367 966 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=144130 $D=1
M312 368 964 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=134870 $D=1
M313 369 965 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=139500 $D=1
M314 370 966 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=144130 $D=1
M315 365 359 368 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=134870 $D=1
M316 366 360 369 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=139500 $D=1
M317 367 361 370 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=144130 $D=1
M318 368 44 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=134870 $D=1
M319 369 44 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=139500 $D=1
M320 370 44 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=144130 $D=1
M321 251 45 368 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=134870 $D=1
M322 252 45 369 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=139500 $D=1
M323 253 45 370 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=144130 $D=1
M324 371 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=134870 $D=1
M325 372 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=139500 $D=1
M326 373 45 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=144130 $D=1
M327 8 46 374 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=134870 $D=1
M328 9 46 375 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=139500 $D=1
M329 140 46 376 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=144130 $D=1
M330 377 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=134870 $D=1
M331 378 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=139500 $D=1
M332 379 47 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=144130 $D=1
M333 380 46 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=134870 $D=1
M334 381 46 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=139500 $D=1
M335 382 46 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=144130 $D=1
M336 8 380 967 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=134870 $D=1
M337 9 381 968 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=139500 $D=1
M338 140 382 969 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=144130 $D=1
M339 383 967 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=134870 $D=1
M340 384 968 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=139500 $D=1
M341 385 969 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=144130 $D=1
M342 380 374 383 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=134870 $D=1
M343 381 375 384 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=139500 $D=1
M344 382 376 385 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=144130 $D=1
M345 383 47 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=134870 $D=1
M346 384 47 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=139500 $D=1
M347 385 47 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=144130 $D=1
M348 251 48 383 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=134870 $D=1
M349 252 48 384 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=139500 $D=1
M350 253 48 385 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=144130 $D=1
M351 386 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=134870 $D=1
M352 387 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=139500 $D=1
M353 388 48 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=144130 $D=1
M354 8 49 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=134870 $D=1
M355 9 49 390 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=139500 $D=1
M356 140 49 391 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=144130 $D=1
M357 392 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=134870 $D=1
M358 393 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=139500 $D=1
M359 394 50 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=144130 $D=1
M360 395 49 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=134870 $D=1
M361 396 49 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=139500 $D=1
M362 397 49 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=144130 $D=1
M363 8 395 970 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=134870 $D=1
M364 9 396 971 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=139500 $D=1
M365 140 397 972 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=144130 $D=1
M366 398 970 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=134870 $D=1
M367 399 971 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=139500 $D=1
M368 400 972 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=144130 $D=1
M369 395 389 398 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=134870 $D=1
M370 396 390 399 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=139500 $D=1
M371 397 391 400 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=144130 $D=1
M372 398 50 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=134870 $D=1
M373 399 50 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=139500 $D=1
M374 400 50 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=144130 $D=1
M375 251 51 398 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=134870 $D=1
M376 252 51 399 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=139500 $D=1
M377 253 51 400 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=144130 $D=1
M378 401 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=134870 $D=1
M379 402 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=139500 $D=1
M380 403 51 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=144130 $D=1
M381 8 52 404 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=134870 $D=1
M382 9 52 405 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=139500 $D=1
M383 140 52 406 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=144130 $D=1
M384 407 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=134870 $D=1
M385 408 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=139500 $D=1
M386 409 53 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=144130 $D=1
M387 410 52 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=134870 $D=1
M388 411 52 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=139500 $D=1
M389 412 52 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=144130 $D=1
M390 8 410 973 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=134870 $D=1
M391 9 411 974 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=139500 $D=1
M392 140 412 975 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=144130 $D=1
M393 413 973 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=134870 $D=1
M394 414 974 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=139500 $D=1
M395 415 975 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=144130 $D=1
M396 410 404 413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=134870 $D=1
M397 411 405 414 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=139500 $D=1
M398 412 406 415 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=144130 $D=1
M399 413 53 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=134870 $D=1
M400 414 53 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=139500 $D=1
M401 415 53 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=144130 $D=1
M402 251 54 413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=134870 $D=1
M403 252 54 414 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=139500 $D=1
M404 253 54 415 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=144130 $D=1
M405 416 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=134870 $D=1
M406 417 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=139500 $D=1
M407 418 54 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=144130 $D=1
M408 8 55 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=134870 $D=1
M409 9 55 420 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=139500 $D=1
M410 140 55 421 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=144130 $D=1
M411 422 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=134870 $D=1
M412 423 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=139500 $D=1
M413 424 56 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=144130 $D=1
M414 425 55 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=134870 $D=1
M415 426 55 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=139500 $D=1
M416 427 55 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=144130 $D=1
M417 8 425 976 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=134870 $D=1
M418 9 426 977 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=139500 $D=1
M419 140 427 978 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=144130 $D=1
M420 428 976 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=134870 $D=1
M421 429 977 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=139500 $D=1
M422 430 978 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=144130 $D=1
M423 425 419 428 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=134870 $D=1
M424 426 420 429 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=139500 $D=1
M425 427 421 430 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=144130 $D=1
M426 428 56 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=134870 $D=1
M427 429 56 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=139500 $D=1
M428 430 56 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=144130 $D=1
M429 251 57 428 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=134870 $D=1
M430 252 57 429 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=139500 $D=1
M431 253 57 430 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=144130 $D=1
M432 431 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=134870 $D=1
M433 432 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=139500 $D=1
M434 433 57 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=144130 $D=1
M435 8 58 434 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=134870 $D=1
M436 9 58 435 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=139500 $D=1
M437 140 58 436 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=144130 $D=1
M438 437 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=134870 $D=1
M439 438 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=139500 $D=1
M440 439 59 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=144130 $D=1
M441 440 58 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=134870 $D=1
M442 441 58 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=139500 $D=1
M443 442 58 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=144130 $D=1
M444 8 440 979 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=134870 $D=1
M445 9 441 980 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=139500 $D=1
M446 140 442 981 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=144130 $D=1
M447 443 979 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=134870 $D=1
M448 444 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=139500 $D=1
M449 445 981 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=144130 $D=1
M450 440 434 443 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=134870 $D=1
M451 441 435 444 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=139500 $D=1
M452 442 436 445 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=144130 $D=1
M453 443 59 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=134870 $D=1
M454 444 59 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=139500 $D=1
M455 445 59 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=144130 $D=1
M456 251 60 443 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=134870 $D=1
M457 252 60 444 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=139500 $D=1
M458 253 60 445 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=144130 $D=1
M459 446 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=134870 $D=1
M460 447 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=139500 $D=1
M461 448 60 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=144130 $D=1
M462 8 61 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=134870 $D=1
M463 9 61 450 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=139500 $D=1
M464 140 61 451 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=144130 $D=1
M465 452 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=134870 $D=1
M466 453 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=139500 $D=1
M467 454 62 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=144130 $D=1
M468 455 61 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=134870 $D=1
M469 456 61 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=139500 $D=1
M470 457 61 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=144130 $D=1
M471 8 455 982 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=134870 $D=1
M472 9 456 983 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=139500 $D=1
M473 140 457 984 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=144130 $D=1
M474 458 982 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=134870 $D=1
M475 459 983 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=139500 $D=1
M476 460 984 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=144130 $D=1
M477 455 449 458 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=134870 $D=1
M478 456 450 459 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=139500 $D=1
M479 457 451 460 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=144130 $D=1
M480 458 62 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=134870 $D=1
M481 459 62 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=139500 $D=1
M482 460 62 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=144130 $D=1
M483 251 63 458 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=134870 $D=1
M484 252 63 459 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=139500 $D=1
M485 253 63 460 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=144130 $D=1
M486 461 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=134870 $D=1
M487 462 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=139500 $D=1
M488 463 63 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=144130 $D=1
M489 8 64 464 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=134870 $D=1
M490 9 64 465 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=139500 $D=1
M491 140 64 466 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=144130 $D=1
M492 467 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=134870 $D=1
M493 468 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=139500 $D=1
M494 469 65 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=144130 $D=1
M495 470 64 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=134870 $D=1
M496 471 64 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=139500 $D=1
M497 472 64 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=144130 $D=1
M498 8 470 985 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=134870 $D=1
M499 9 471 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=139500 $D=1
M500 140 472 987 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=144130 $D=1
M501 473 985 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=134870 $D=1
M502 474 986 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=139500 $D=1
M503 475 987 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=144130 $D=1
M504 470 464 473 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=134870 $D=1
M505 471 465 474 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=139500 $D=1
M506 472 466 475 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=144130 $D=1
M507 473 65 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=134870 $D=1
M508 474 65 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=139500 $D=1
M509 475 65 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=144130 $D=1
M510 251 66 473 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=134870 $D=1
M511 252 66 474 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=139500 $D=1
M512 253 66 475 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=144130 $D=1
M513 476 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=134870 $D=1
M514 477 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=139500 $D=1
M515 478 66 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=144130 $D=1
M516 8 67 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=134870 $D=1
M517 9 67 480 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=139500 $D=1
M518 140 67 481 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=144130 $D=1
M519 482 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=134870 $D=1
M520 483 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=139500 $D=1
M521 484 68 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=144130 $D=1
M522 485 67 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=134870 $D=1
M523 486 67 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=139500 $D=1
M524 487 67 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=144130 $D=1
M525 8 485 988 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=134870 $D=1
M526 9 486 989 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=139500 $D=1
M527 140 487 990 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=144130 $D=1
M528 488 988 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=134870 $D=1
M529 489 989 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=139500 $D=1
M530 490 990 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=144130 $D=1
M531 485 479 488 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=134870 $D=1
M532 486 480 489 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=139500 $D=1
M533 487 481 490 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=144130 $D=1
M534 488 68 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=134870 $D=1
M535 489 68 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=139500 $D=1
M536 490 68 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=144130 $D=1
M537 251 69 488 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=134870 $D=1
M538 252 69 489 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=139500 $D=1
M539 253 69 490 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=144130 $D=1
M540 491 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=134870 $D=1
M541 492 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=139500 $D=1
M542 493 69 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=144130 $D=1
M543 8 70 494 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=134870 $D=1
M544 9 70 495 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=139500 $D=1
M545 140 70 496 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=144130 $D=1
M546 497 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=134870 $D=1
M547 498 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=139500 $D=1
M548 499 71 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=144130 $D=1
M549 500 70 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=134870 $D=1
M550 501 70 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=139500 $D=1
M551 502 70 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=144130 $D=1
M552 8 500 991 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=134870 $D=1
M553 9 501 992 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=139500 $D=1
M554 140 502 993 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=144130 $D=1
M555 503 991 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=134870 $D=1
M556 504 992 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=139500 $D=1
M557 505 993 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=144130 $D=1
M558 500 494 503 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=134870 $D=1
M559 501 495 504 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=139500 $D=1
M560 502 496 505 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=144130 $D=1
M561 503 71 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=134870 $D=1
M562 504 71 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=139500 $D=1
M563 505 71 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=144130 $D=1
M564 251 72 503 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=134870 $D=1
M565 252 72 504 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=139500 $D=1
M566 253 72 505 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=144130 $D=1
M567 506 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=134870 $D=1
M568 507 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=139500 $D=1
M569 508 72 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=144130 $D=1
M570 8 73 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=134870 $D=1
M571 9 73 510 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=139500 $D=1
M572 140 73 511 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=144130 $D=1
M573 512 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=134870 $D=1
M574 513 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=139500 $D=1
M575 514 74 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=144130 $D=1
M576 515 73 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=134870 $D=1
M577 516 73 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=139500 $D=1
M578 517 73 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=144130 $D=1
M579 8 515 994 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=134870 $D=1
M580 9 516 995 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=139500 $D=1
M581 140 517 996 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=144130 $D=1
M582 518 994 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=134870 $D=1
M583 519 995 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=139500 $D=1
M584 520 996 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=144130 $D=1
M585 515 509 518 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=134870 $D=1
M586 516 510 519 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=139500 $D=1
M587 517 511 520 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=144130 $D=1
M588 518 74 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=134870 $D=1
M589 519 74 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=139500 $D=1
M590 520 74 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=144130 $D=1
M591 251 75 518 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=134870 $D=1
M592 252 75 519 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=139500 $D=1
M593 253 75 520 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=144130 $D=1
M594 521 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=134870 $D=1
M595 522 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=139500 $D=1
M596 523 75 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=144130 $D=1
M597 8 76 524 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=134870 $D=1
M598 9 76 525 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=139500 $D=1
M599 140 76 526 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=144130 $D=1
M600 527 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=134870 $D=1
M601 528 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=139500 $D=1
M602 529 77 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=144130 $D=1
M603 530 76 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=134870 $D=1
M604 531 76 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=139500 $D=1
M605 532 76 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=144130 $D=1
M606 8 530 997 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=134870 $D=1
M607 9 531 998 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=139500 $D=1
M608 140 532 999 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=144130 $D=1
M609 533 997 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=134870 $D=1
M610 534 998 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=139500 $D=1
M611 535 999 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=144130 $D=1
M612 530 524 533 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=134870 $D=1
M613 531 525 534 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=139500 $D=1
M614 532 526 535 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=144130 $D=1
M615 533 77 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=134870 $D=1
M616 534 77 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=139500 $D=1
M617 535 77 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=144130 $D=1
M618 251 78 533 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=134870 $D=1
M619 252 78 534 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=139500 $D=1
M620 253 78 535 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=144130 $D=1
M621 536 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=134870 $D=1
M622 537 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=139500 $D=1
M623 538 78 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=144130 $D=1
M624 8 79 539 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=134870 $D=1
M625 9 79 540 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=139500 $D=1
M626 140 79 541 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=144130 $D=1
M627 542 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=134870 $D=1
M628 543 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=139500 $D=1
M629 544 80 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=144130 $D=1
M630 545 79 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=134870 $D=1
M631 546 79 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=139500 $D=1
M632 547 79 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=144130 $D=1
M633 8 545 1000 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=134870 $D=1
M634 9 546 1001 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=139500 $D=1
M635 140 547 1002 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=144130 $D=1
M636 548 1000 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=134870 $D=1
M637 549 1001 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=139500 $D=1
M638 550 1002 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=144130 $D=1
M639 545 539 548 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=134870 $D=1
M640 546 540 549 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=139500 $D=1
M641 547 541 550 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=144130 $D=1
M642 548 80 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=134870 $D=1
M643 549 80 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=139500 $D=1
M644 550 80 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=144130 $D=1
M645 251 81 548 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=134870 $D=1
M646 252 81 549 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=139500 $D=1
M647 253 81 550 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=144130 $D=1
M648 551 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=134870 $D=1
M649 552 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=139500 $D=1
M650 553 81 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=144130 $D=1
M651 8 82 554 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=134870 $D=1
M652 9 82 555 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=139500 $D=1
M653 140 82 556 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=144130 $D=1
M654 557 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=134870 $D=1
M655 558 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=139500 $D=1
M656 559 83 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=144130 $D=1
M657 560 82 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=134870 $D=1
M658 561 82 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=139500 $D=1
M659 562 82 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=144130 $D=1
M660 8 560 1003 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=134870 $D=1
M661 9 561 1004 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=139500 $D=1
M662 140 562 1005 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=144130 $D=1
M663 563 1003 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=134870 $D=1
M664 564 1004 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=139500 $D=1
M665 565 1005 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=144130 $D=1
M666 560 554 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=134870 $D=1
M667 561 555 564 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=139500 $D=1
M668 562 556 565 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=144130 $D=1
M669 563 83 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=134870 $D=1
M670 564 83 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=139500 $D=1
M671 565 83 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=144130 $D=1
M672 251 84 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=134870 $D=1
M673 252 84 564 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=139500 $D=1
M674 253 84 565 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=144130 $D=1
M675 566 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=134870 $D=1
M676 567 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=139500 $D=1
M677 568 84 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=144130 $D=1
M678 8 85 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=134870 $D=1
M679 9 85 570 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=139500 $D=1
M680 140 85 571 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=144130 $D=1
M681 572 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=134870 $D=1
M682 573 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=139500 $D=1
M683 574 86 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=144130 $D=1
M684 575 85 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=134870 $D=1
M685 576 85 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=139500 $D=1
M686 577 85 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=144130 $D=1
M687 8 575 1006 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=134870 $D=1
M688 9 576 1007 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=139500 $D=1
M689 140 577 1008 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=144130 $D=1
M690 578 1006 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=134870 $D=1
M691 579 1007 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=139500 $D=1
M692 580 1008 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=144130 $D=1
M693 575 569 578 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=134870 $D=1
M694 576 570 579 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=139500 $D=1
M695 577 571 580 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=144130 $D=1
M696 578 86 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=134870 $D=1
M697 579 86 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=139500 $D=1
M698 580 86 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=144130 $D=1
M699 251 87 578 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=134870 $D=1
M700 252 87 579 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=139500 $D=1
M701 253 87 580 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=144130 $D=1
M702 581 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=134870 $D=1
M703 582 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=139500 $D=1
M704 583 87 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=144130 $D=1
M705 8 88 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=134870 $D=1
M706 9 88 585 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=139500 $D=1
M707 140 88 586 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=144130 $D=1
M708 587 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=134870 $D=1
M709 588 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=139500 $D=1
M710 589 89 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=144130 $D=1
M711 590 88 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=134870 $D=1
M712 591 88 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=139500 $D=1
M713 592 88 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=144130 $D=1
M714 8 590 1009 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=134870 $D=1
M715 9 591 1010 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=139500 $D=1
M716 140 592 1011 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=144130 $D=1
M717 593 1009 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=134870 $D=1
M718 594 1010 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=139500 $D=1
M719 595 1011 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=144130 $D=1
M720 590 584 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=134870 $D=1
M721 591 585 594 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=139500 $D=1
M722 592 586 595 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=144130 $D=1
M723 593 89 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=134870 $D=1
M724 594 89 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=139500 $D=1
M725 595 89 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=144130 $D=1
M726 251 90 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=134870 $D=1
M727 252 90 594 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=139500 $D=1
M728 253 90 595 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=144130 $D=1
M729 596 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=134870 $D=1
M730 597 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=139500 $D=1
M731 598 90 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=144130 $D=1
M732 8 91 599 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=134870 $D=1
M733 9 91 600 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=139500 $D=1
M734 140 91 601 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=144130 $D=1
M735 602 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=134870 $D=1
M736 603 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=139500 $D=1
M737 604 92 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=144130 $D=1
M738 605 91 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=134870 $D=1
M739 606 91 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=139500 $D=1
M740 607 91 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=144130 $D=1
M741 8 605 1012 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=134870 $D=1
M742 9 606 1013 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=139500 $D=1
M743 140 607 1014 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=144130 $D=1
M744 608 1012 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=134870 $D=1
M745 609 1013 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=139500 $D=1
M746 610 1014 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=144130 $D=1
M747 605 599 608 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=134870 $D=1
M748 606 600 609 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=139500 $D=1
M749 607 601 610 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=144130 $D=1
M750 608 92 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=134870 $D=1
M751 609 92 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=139500 $D=1
M752 610 92 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=144130 $D=1
M753 251 93 608 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=134870 $D=1
M754 252 93 609 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=139500 $D=1
M755 253 93 610 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=144130 $D=1
M756 611 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=134870 $D=1
M757 612 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=139500 $D=1
M758 613 93 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=144130 $D=1
M759 8 94 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=134870 $D=1
M760 9 94 615 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=139500 $D=1
M761 140 94 616 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=144130 $D=1
M762 617 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=134870 $D=1
M763 618 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=139500 $D=1
M764 619 95 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=144130 $D=1
M765 620 94 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=134870 $D=1
M766 621 94 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=139500 $D=1
M767 622 94 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=144130 $D=1
M768 8 620 1015 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=134870 $D=1
M769 9 621 1016 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=139500 $D=1
M770 140 622 1017 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=144130 $D=1
M771 623 1015 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=134870 $D=1
M772 624 1016 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=139500 $D=1
M773 625 1017 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=144130 $D=1
M774 620 614 623 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=134870 $D=1
M775 621 615 624 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=139500 $D=1
M776 622 616 625 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=144130 $D=1
M777 623 95 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=134870 $D=1
M778 624 95 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=139500 $D=1
M779 625 95 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=144130 $D=1
M780 251 96 623 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=134870 $D=1
M781 252 96 624 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=139500 $D=1
M782 253 96 625 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=144130 $D=1
M783 626 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=134870 $D=1
M784 627 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=139500 $D=1
M785 628 96 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=144130 $D=1
M786 8 97 629 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=134870 $D=1
M787 9 97 630 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=139500 $D=1
M788 140 97 631 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=144130 $D=1
M789 632 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=134870 $D=1
M790 633 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=139500 $D=1
M791 634 98 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=144130 $D=1
M792 635 97 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=134870 $D=1
M793 636 97 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=139500 $D=1
M794 637 97 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=144130 $D=1
M795 8 635 1018 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=134870 $D=1
M796 9 636 1019 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=139500 $D=1
M797 140 637 1020 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=144130 $D=1
M798 638 1018 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=134870 $D=1
M799 639 1019 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=139500 $D=1
M800 640 1020 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=144130 $D=1
M801 635 629 638 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=134870 $D=1
M802 636 630 639 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=139500 $D=1
M803 637 631 640 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=144130 $D=1
M804 638 98 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=134870 $D=1
M805 639 98 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=139500 $D=1
M806 640 98 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=144130 $D=1
M807 251 99 638 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=134870 $D=1
M808 252 99 639 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=139500 $D=1
M809 253 99 640 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=144130 $D=1
M810 641 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=134870 $D=1
M811 642 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=139500 $D=1
M812 643 99 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=144130 $D=1
M813 8 100 644 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=134870 $D=1
M814 9 100 645 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=139500 $D=1
M815 140 100 646 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=144130 $D=1
M816 647 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=134870 $D=1
M817 648 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=139500 $D=1
M818 649 101 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=144130 $D=1
M819 650 100 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=134870 $D=1
M820 651 100 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=139500 $D=1
M821 652 100 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=144130 $D=1
M822 8 650 1021 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=134870 $D=1
M823 9 651 1022 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=139500 $D=1
M824 140 652 1023 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=144130 $D=1
M825 653 1021 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=134870 $D=1
M826 654 1022 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=139500 $D=1
M827 655 1023 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=144130 $D=1
M828 650 644 653 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=134870 $D=1
M829 651 645 654 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=139500 $D=1
M830 652 646 655 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=144130 $D=1
M831 653 101 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=134870 $D=1
M832 654 101 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=139500 $D=1
M833 655 101 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=144130 $D=1
M834 251 102 653 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=134870 $D=1
M835 252 102 654 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=139500 $D=1
M836 253 102 655 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=144130 $D=1
M837 656 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=134870 $D=1
M838 657 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=139500 $D=1
M839 658 102 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=144130 $D=1
M840 8 103 659 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=134870 $D=1
M841 9 103 660 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=139500 $D=1
M842 140 103 661 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=144130 $D=1
M843 662 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=134870 $D=1
M844 663 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=139500 $D=1
M845 664 104 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=144130 $D=1
M846 665 103 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=134870 $D=1
M847 666 103 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=139500 $D=1
M848 667 103 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=144130 $D=1
M849 8 665 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=134870 $D=1
M850 9 666 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=139500 $D=1
M851 140 667 1026 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=144130 $D=1
M852 668 1024 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=134870 $D=1
M853 669 1025 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=139500 $D=1
M854 670 1026 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=144130 $D=1
M855 665 659 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=134870 $D=1
M856 666 660 669 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=139500 $D=1
M857 667 661 670 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=144130 $D=1
M858 668 104 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=134870 $D=1
M859 669 104 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=139500 $D=1
M860 670 104 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=144130 $D=1
M861 251 105 668 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=134870 $D=1
M862 252 105 669 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=139500 $D=1
M863 253 105 670 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=144130 $D=1
M864 671 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=134870 $D=1
M865 672 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=139500 $D=1
M866 673 105 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=144130 $D=1
M867 8 106 674 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=134870 $D=1
M868 9 106 675 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=139500 $D=1
M869 140 106 676 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=144130 $D=1
M870 677 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=134870 $D=1
M871 678 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=139500 $D=1
M872 679 107 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=144130 $D=1
M873 680 106 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=134870 $D=1
M874 681 106 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=139500 $D=1
M875 682 106 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=144130 $D=1
M876 8 680 1027 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=134870 $D=1
M877 9 681 1028 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=139500 $D=1
M878 140 682 1029 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=144130 $D=1
M879 683 1027 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=134870 $D=1
M880 684 1028 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=139500 $D=1
M881 685 1029 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=144130 $D=1
M882 680 674 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=134870 $D=1
M883 681 675 684 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=139500 $D=1
M884 682 676 685 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=144130 $D=1
M885 683 107 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=134870 $D=1
M886 684 107 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=139500 $D=1
M887 685 107 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=144130 $D=1
M888 251 108 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=134870 $D=1
M889 252 108 684 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=139500 $D=1
M890 253 108 685 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=144130 $D=1
M891 686 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=134870 $D=1
M892 687 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=139500 $D=1
M893 688 108 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=144130 $D=1
M894 8 109 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=134870 $D=1
M895 9 109 690 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=139500 $D=1
M896 140 109 691 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=144130 $D=1
M897 692 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=134870 $D=1
M898 693 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=139500 $D=1
M899 694 110 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=144130 $D=1
M900 695 109 230 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=134870 $D=1
M901 696 109 231 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=139500 $D=1
M902 697 109 232 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=144130 $D=1
M903 8 695 1030 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=134870 $D=1
M904 9 696 1031 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=139500 $D=1
M905 140 697 1032 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=144130 $D=1
M906 698 1030 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=134870 $D=1
M907 699 1031 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=139500 $D=1
M908 700 1032 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=144130 $D=1
M909 695 689 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=134870 $D=1
M910 696 690 699 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=139500 $D=1
M911 697 691 700 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=144130 $D=1
M912 698 110 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=134870 $D=1
M913 699 110 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=139500 $D=1
M914 700 110 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=144130 $D=1
M915 251 111 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=134870 $D=1
M916 252 111 699 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=139500 $D=1
M917 253 111 700 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=144130 $D=1
M918 701 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=134870 $D=1
M919 702 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=139500 $D=1
M920 703 111 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=144130 $D=1
M921 8 112 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=134870 $D=1
M922 9 112 705 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=139500 $D=1
M923 140 112 706 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=144130 $D=1
M924 707 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=134870 $D=1
M925 708 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=139500 $D=1
M926 709 113 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=144130 $D=1
M927 8 113 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=134870 $D=1
M928 9 113 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=139500 $D=1
M929 140 113 247 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=144130 $D=1
M930 251 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=134870 $D=1
M931 252 112 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=139500 $D=1
M932 253 112 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=144130 $D=1
M933 8 713 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=134870 $D=1
M934 9 714 711 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=139500 $D=1
M935 140 715 712 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=144130 $D=1
M936 713 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=134870 $D=1
M937 714 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=139500 $D=1
M938 715 114 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=144130 $D=1
M939 1033 245 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=134870 $D=1
M940 1034 246 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=139500 $D=1
M941 1035 247 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=144130 $D=1
M942 716 710 1033 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=134870 $D=1
M943 717 711 1034 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=139500 $D=1
M944 718 712 1035 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=144130 $D=1
M945 8 716 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=134870 $D=1
M946 9 717 720 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=139500 $D=1
M947 140 718 721 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=144130 $D=1
M948 1036 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=134870 $D=1
M949 1037 720 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=139500 $D=1
M950 1038 721 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=144130 $D=1
M951 716 713 1036 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=134870 $D=1
M952 717 714 1037 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=139500 $D=1
M953 718 715 1038 140 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=144130 $D=1
M954 8 725 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=134870 $D=1
M955 9 726 723 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=139500 $D=1
M956 140 727 724 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=144130 $D=1
M957 725 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=134870 $D=1
M958 726 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=139500 $D=1
M959 727 114 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=144130 $D=1
M960 1039 251 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=134870 $D=1
M961 1040 252 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=139500 $D=1
M962 1041 253 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=144130 $D=1
M963 728 722 1039 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=134870 $D=1
M964 729 723 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=139500 $D=1
M965 730 724 1041 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=144130 $D=1
M966 8 728 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=134870 $D=1
M967 9 729 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=139500 $D=1
M968 140 730 117 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=144130 $D=1
M969 1042 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=134870 $D=1
M970 1043 116 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=139500 $D=1
M971 1044 117 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=144130 $D=1
M972 728 725 1042 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=134870 $D=1
M973 729 726 1043 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=139500 $D=1
M974 730 727 1044 140 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=144130 $D=1
M975 731 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=134870 $D=1
M976 732 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=139500 $D=1
M977 733 118 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=144130 $D=1
M978 734 731 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=134870 $D=1
M979 735 732 720 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=139500 $D=1
M980 736 733 721 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=144130 $D=1
M981 119 118 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=134870 $D=1
M982 120 118 735 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=139500 $D=1
M983 121 118 736 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=144130 $D=1
M984 737 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=134870 $D=1
M985 738 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=139500 $D=1
M986 739 122 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=144130 $D=1
M987 740 737 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=134870 $D=1
M988 741 738 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=139500 $D=1
M989 742 739 117 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=144130 $D=1
M990 1045 122 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=134870 $D=1
M991 1046 122 741 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=139500 $D=1
M992 1047 122 742 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=144130 $D=1
M993 8 115 1045 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=134870 $D=1
M994 9 116 1046 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=139500 $D=1
M995 140 117 1047 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=144130 $D=1
M996 743 123 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=134870 $D=1
M997 744 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=139500 $D=1
M998 745 123 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=144130 $D=1
M999 124 743 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=134870 $D=1
M1000 125 744 741 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=139500 $D=1
M1001 126 745 742 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=144130 $D=1
M1002 11 123 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=134870 $D=1
M1003 12 123 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=139500 $D=1
M1004 13 123 126 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=144130 $D=1
M1005 748 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=134870 $D=1
M1006 749 747 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=139500 $D=1
M1007 750 127 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=144130 $D=1
M1008 8 754 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=134870 $D=1
M1009 9 755 752 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=139500 $D=1
M1010 140 756 753 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=144130 $D=1
M1011 757 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=134870 $D=1
M1012 758 735 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=139500 $D=1
M1013 759 736 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=144130 $D=1
M1014 754 757 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=134870 $D=1
M1015 755 758 747 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=139500 $D=1
M1016 756 759 127 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=144130 $D=1
M1017 748 734 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=134870 $D=1
M1018 749 735 755 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=139500 $D=1
M1019 750 736 756 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=144130 $D=1
M1020 760 751 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=134870 $D=1
M1021 761 752 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=139500 $D=1
M1022 762 753 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=144130 $D=1
M1023 128 760 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=134870 $D=1
M1024 746 761 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=139500 $D=1
M1025 747 762 126 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=144130 $D=1
M1026 734 751 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=134870 $D=1
M1027 735 752 746 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=139500 $D=1
M1028 736 753 747 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=144130 $D=1
M1029 763 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=134870 $D=1
M1030 764 746 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=139500 $D=1
M1031 765 747 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=144130 $D=1
M1032 766 751 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=134870 $D=1
M1033 767 752 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=139500 $D=1
M1034 768 753 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=144130 $D=1
M1035 769 766 763 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=134870 $D=1
M1036 770 767 764 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=139500 $D=1
M1037 771 768 765 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=144130 $D=1
M1038 124 751 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=134870 $D=1
M1039 125 752 770 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=139500 $D=1
M1040 126 753 771 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=144130 $D=1
M1041 772 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=134870 $D=1
M1042 773 735 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=139500 $D=1
M1043 774 736 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=144130 $D=1
M1044 8 124 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=134870 $D=1
M1045 9 125 773 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=139500 $D=1
M1046 140 126 774 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=144130 $D=1
M1047 775 769 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=134870 $D=1
M1048 776 770 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=139500 $D=1
M1049 777 771 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=144130 $D=1
M1050 1075 734 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=134870 $D=1
M1051 1076 735 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=139500 $D=1
M1052 1077 736 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=144130 $D=1
M1053 778 124 1075 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=134870 $D=1
M1054 779 125 1076 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=139500 $D=1
M1055 780 126 1077 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=144130 $D=1
M1056 1078 734 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=134870 $D=1
M1057 1079 735 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=139500 $D=1
M1058 1080 736 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=144130 $D=1
M1059 781 124 1078 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=134870 $D=1
M1060 782 125 1079 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=139500 $D=1
M1061 783 126 1080 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=144130 $D=1
M1062 787 734 784 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=134870 $D=1
M1063 788 735 785 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=139500 $D=1
M1064 789 736 786 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=144130 $D=1
M1065 784 124 787 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=134870 $D=1
M1066 785 125 788 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=139500 $D=1
M1067 786 126 789 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=144130 $D=1
M1068 8 781 784 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=134870 $D=1
M1069 9 782 785 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=139500 $D=1
M1070 140 783 786 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=144130 $D=1
M1071 790 135 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=134870 $D=1
M1072 791 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=139500 $D=1
M1073 792 135 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=144130 $D=1
M1074 793 790 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=134870 $D=1
M1075 794 791 773 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=139500 $D=1
M1076 795 792 774 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=144130 $D=1
M1077 778 135 793 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=134870 $D=1
M1078 779 135 794 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=139500 $D=1
M1079 780 135 795 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=144130 $D=1
M1080 796 790 775 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=134870 $D=1
M1081 797 791 776 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=139500 $D=1
M1082 798 792 777 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=144130 $D=1
M1083 787 135 796 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=134870 $D=1
M1084 788 135 797 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=139500 $D=1
M1085 789 135 798 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=144130 $D=1
M1086 799 136 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=134870 $D=1
M1087 800 136 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=139500 $D=1
M1088 801 136 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=144130 $D=1
M1089 802 799 796 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=134870 $D=1
M1090 803 800 797 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=139500 $D=1
M1091 804 801 798 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=144130 $D=1
M1092 793 136 802 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=134870 $D=1
M1093 794 136 803 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=139500 $D=1
M1094 795 136 804 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=144130 $D=1
M1095 14 802 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=134870 $D=1
M1096 15 803 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=139500 $D=1
M1097 16 804 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=144130 $D=1
M1098 805 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=134870 $D=1
M1099 806 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=139500 $D=1
M1100 807 137 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=144130 $D=1
M1101 808 805 138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=134870 $D=1
M1102 809 806 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=139500 $D=1
M1103 810 807 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=144130 $D=1
M1104 141 137 808 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=134870 $D=1
M1105 142 137 809 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=139500 $D=1
M1106 138 137 810 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=144130 $D=1
M1107 811 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=134870 $D=1
M1108 812 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=139500 $D=1
M1109 813 137 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=144130 $D=1
M1110 814 811 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=134870 $D=1
M1111 815 812 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=139500 $D=1
M1112 816 813 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=144130 $D=1
M1113 144 137 814 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=134870 $D=1
M1114 145 137 815 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=139500 $D=1
M1115 146 137 816 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=144130 $D=1
M1116 817 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=134870 $D=1
M1117 818 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=139500 $D=1
M1118 819 137 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=144130 $D=1
M1119 820 817 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=134870 $D=1
M1120 821 818 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=139500 $D=1
M1121 822 819 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=144130 $D=1
M1122 147 137 820 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=134870 $D=1
M1123 148 137 821 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=139500 $D=1
M1124 149 137 822 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=144130 $D=1
M1125 823 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=134870 $D=1
M1126 824 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=139500 $D=1
M1127 825 137 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=144130 $D=1
M1128 826 823 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=134870 $D=1
M1129 827 824 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=139500 $D=1
M1130 828 825 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=144130 $D=1
M1131 150 137 826 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=134870 $D=1
M1132 151 137 827 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=139500 $D=1
M1133 152 137 828 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=144130 $D=1
M1134 829 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=134870 $D=1
M1135 830 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=139500 $D=1
M1136 831 137 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=144130 $D=1
M1137 832 829 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=134870 $D=1
M1138 833 830 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=139500 $D=1
M1139 834 831 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=144130 $D=1
M1140 153 137 832 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=134870 $D=1
M1141 154 137 833 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=139500 $D=1
M1142 155 137 834 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=144130 $D=1
M1143 8 734 1048 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=134870 $D=1
M1144 9 735 1049 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=139500 $D=1
M1145 140 736 1050 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=144130 $D=1
M1146 142 1048 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=134870 $D=1
M1147 138 1049 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=139500 $D=1
M1148 139 1050 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=144130 $D=1
M1149 835 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=134870 $D=1
M1150 836 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=139500 $D=1
M1151 837 126 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=144130 $D=1
M1152 146 835 142 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=134870 $D=1
M1153 156 836 138 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=139500 $D=1
M1154 143 837 139 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=144130 $D=1
M1155 808 126 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=134870 $D=1
M1156 809 126 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=139500 $D=1
M1157 810 126 143 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=144130 $D=1
M1158 838 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=134870 $D=1
M1159 839 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=139500 $D=1
M1160 840 125 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=144130 $D=1
M1161 134 838 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=134870 $D=1
M1162 133 839 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=139500 $D=1
M1163 132 840 143 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=144130 $D=1
M1164 814 125 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=134870 $D=1
M1165 815 125 133 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=139500 $D=1
M1166 816 125 132 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=144130 $D=1
M1167 841 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=134870 $D=1
M1168 842 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=139500 $D=1
M1169 843 124 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=144130 $D=1
M1170 129 841 134 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=134870 $D=1
M1171 130 842 133 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=139500 $D=1
M1172 131 843 132 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=144130 $D=1
M1173 820 124 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=134870 $D=1
M1174 821 124 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=139500 $D=1
M1175 822 124 131 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=144130 $D=1
M1176 844 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=134870 $D=1
M1177 845 157 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=139500 $D=1
M1178 846 157 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=144130 $D=1
M1179 158 844 129 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=134870 $D=1
M1180 159 845 130 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=139500 $D=1
M1181 160 846 131 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=144130 $D=1
M1182 826 157 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=134870 $D=1
M1183 827 157 159 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=139500 $D=1
M1184 828 157 160 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=144130 $D=1
M1185 847 161 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=134870 $D=1
M1186 848 161 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=139500 $D=1
M1187 849 161 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=144130 $D=1
M1188 209 847 158 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=134870 $D=1
M1189 210 848 159 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=139500 $D=1
M1190 211 849 160 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=144130 $D=1
M1191 832 161 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=134870 $D=1
M1192 833 161 210 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=139500 $D=1
M1193 834 161 211 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=144130 $D=1
M1194 850 162 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=134870 $D=1
M1195 851 162 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=139500 $D=1
M1196 852 162 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=144130 $D=1
M1197 853 850 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=134870 $D=1
M1198 854 851 116 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=139500 $D=1
M1199 855 852 117 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=144130 $D=1
M1200 11 162 853 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=134870 $D=1
M1201 12 162 854 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=139500 $D=1
M1202 13 162 855 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=144130 $D=1
M1203 1081 719 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=134870 $D=1
M1204 1082 720 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=139500 $D=1
M1205 1083 721 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=144130 $D=1
M1206 856 853 1081 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=134870 $D=1
M1207 857 854 1082 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=139500 $D=1
M1208 858 855 1083 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=144130 $D=1
M1209 862 719 859 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=134870 $D=1
M1210 863 720 860 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=139500 $D=1
M1211 864 721 861 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=144130 $D=1
M1212 859 853 862 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=134870 $D=1
M1213 860 854 863 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=139500 $D=1
M1214 861 855 864 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=144130 $D=1
M1215 8 856 859 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=134870 $D=1
M1216 9 857 860 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=139500 $D=1
M1217 140 858 861 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=144130 $D=1
M1218 1084 163 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=134870 $D=1
M1219 1085 865 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=139500 $D=1
M1220 1086 866 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=144130 $D=1
M1221 1051 862 1084 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=134870 $D=1
M1222 1052 863 1085 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=139500 $D=1
M1223 1053 864 1086 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=144130 $D=1
M1224 865 1051 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=134870 $D=1
M1225 866 1052 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=139500 $D=1
M1226 164 1053 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=144130 $D=1
M1227 867 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=134870 $D=1
M1228 868 720 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=139500 $D=1
M1229 869 721 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=144130 $D=1
M1230 8 870 867 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=134870 $D=1
M1231 9 871 868 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=139500 $D=1
M1232 140 872 869 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=144130 $D=1
M1233 870 853 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=134870 $D=1
M1234 871 854 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=139500 $D=1
M1235 872 855 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=144130 $D=1
M1236 1087 867 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=134870 $D=1
M1237 1088 868 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=139500 $D=1
M1238 1089 869 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=144130 $D=1
M1239 873 163 1087 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=134870 $D=1
M1240 874 865 1088 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=139500 $D=1
M1241 875 866 1089 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=144130 $D=1
M1242 878 165 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=134870 $D=1
M1243 879 876 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=139500 $D=1
M1244 880 877 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=144130 $D=1
M1245 1090 873 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=134870 $D=1
M1246 1091 874 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=139500 $D=1
M1247 1092 875 140 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=144130 $D=1
M1248 876 878 1090 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=134870 $D=1
M1249 877 879 1091 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=139500 $D=1
M1250 166 880 1092 140 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=144130 $D=1
M1251 883 881 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=134870 $D=1
M1252 884 882 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=139500 $D=1
M1253 885 140 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=144130 $D=1
M1254 8 889 886 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=134870 $D=1
M1255 9 890 887 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=139500 $D=1
M1256 140 891 888 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=144130 $D=1
M1257 892 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=134870 $D=1
M1258 893 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=139500 $D=1
M1259 894 121 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=144130 $D=1
M1260 889 892 881 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=134870 $D=1
M1261 890 893 882 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=139500 $D=1
M1262 891 894 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=144130 $D=1
M1263 883 119 889 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=134870 $D=1
M1264 884 120 890 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=139500 $D=1
M1265 885 121 891 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=144130 $D=1
M1266 895 886 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=134870 $D=1
M1267 896 887 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=139500 $D=1
M1268 897 888 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=144130 $D=1
M1269 168 895 167 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=134870 $D=1
M1270 881 896 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=139500 $D=1
M1271 882 897 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=144130 $D=1
M1272 119 886 168 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=134870 $D=1
M1273 120 887 881 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=139500 $D=1
M1274 121 888 882 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=144130 $D=1
M1275 898 168 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=134870 $D=1
M1276 899 881 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=139500 $D=1
M1277 900 882 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=144130 $D=1
M1278 901 886 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=134870 $D=1
M1279 902 887 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=139500 $D=1
M1280 903 888 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=144130 $D=1
M1281 212 901 898 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=134870 $D=1
M1282 213 902 899 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=139500 $D=1
M1283 214 903 900 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=144130 $D=1
M1284 167 886 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=134870 $D=1
M1285 9 887 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=139500 $D=1
M1286 140 888 214 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=144130 $D=1
M1287 904 169 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=134870 $D=1
M1288 905 169 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=139500 $D=1
M1289 906 169 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=144130 $D=1
M1290 907 904 212 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=134870 $D=1
M1291 908 905 213 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=139500 $D=1
M1292 909 906 214 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=144130 $D=1
M1293 14 169 907 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=134870 $D=1
M1294 15 169 908 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=139500 $D=1
M1295 16 169 909 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=144130 $D=1
M1296 910 170 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=134870 $D=1
M1297 911 170 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=139500 $D=1
M1298 912 170 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=144130 $D=1
M1299 170 910 907 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=134870 $D=1
M1300 170 911 908 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=139500 $D=1
M1301 170 912 909 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=144130 $D=1
M1302 8 170 170 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=134870 $D=1
M1303 9 170 170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=139500 $D=1
M1304 140 170 170 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=144130 $D=1
M1305 913 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=134870 $D=1
M1306 914 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=139500 $D=1
M1307 915 114 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=144130 $D=1
M1308 8 913 916 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=134870 $D=1
M1309 9 914 917 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=139500 $D=1
M1310 140 915 918 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=144130 $D=1
M1311 919 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=134870 $D=1
M1312 920 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=139500 $D=1
M1313 921 114 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=144130 $D=1
M1314 922 913 170 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=134870 $D=1
M1315 923 914 170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=139500 $D=1
M1316 924 915 170 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=144130 $D=1
M1317 8 922 1054 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=134870 $D=1
M1318 9 923 1055 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=139500 $D=1
M1319 140 924 1056 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=144130 $D=1
M1320 925 1054 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=134870 $D=1
M1321 926 1055 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=139500 $D=1
M1322 927 1056 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=144130 $D=1
M1323 922 916 925 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=134870 $D=1
M1324 923 917 926 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=139500 $D=1
M1325 924 918 927 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=144130 $D=1
M1326 928 114 925 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=134870 $D=1
M1327 929 114 926 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=139500 $D=1
M1328 930 114 927 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=144130 $D=1
M1329 8 934 931 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=134870 $D=1
M1330 9 935 932 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=139500 $D=1
M1331 140 936 933 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=144130 $D=1
M1332 934 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=134870 $D=1
M1333 935 114 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=139500 $D=1
M1334 936 114 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=144130 $D=1
M1335 1057 928 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=134870 $D=1
M1336 1058 929 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=139500 $D=1
M1337 1059 930 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=144130 $D=1
M1338 937 931 1057 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=134870 $D=1
M1339 938 932 1058 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=139500 $D=1
M1340 939 933 1059 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=144130 $D=1
M1341 8 937 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=134870 $D=1
M1342 9 938 120 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=139500 $D=1
M1343 140 939 121 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=144130 $D=1
M1344 1060 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=134870 $D=1
M1345 1061 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=139500 $D=1
M1346 1062 121 140 140 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=144130 $D=1
M1347 937 934 1060 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=134870 $D=1
M1348 938 935 1061 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=139500 $D=1
M1349 939 936 1062 140 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=144130 $D=1
M1350 173 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=136120 $D=0
M1351 174 1 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=140750 $D=0
M1352 175 1 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=145380 $D=0
M1353 176 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=136120 $D=0
M1354 177 1 3 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=140750 $D=0
M1355 178 1 4 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=145380 $D=0
M1356 8 173 176 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=136120 $D=0
M1357 9 174 177 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=140750 $D=0
M1358 140 175 178 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=145380 $D=0
M1359 179 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=136120 $D=0
M1360 180 1 3 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=140750 $D=0
M1361 181 1 4 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=145380 $D=0
M1362 2 173 179 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=136120 $D=0
M1363 3 174 180 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=140750 $D=0
M1364 4 175 181 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=145380 $D=0
M1365 182 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=136120 $D=0
M1366 183 1 3 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=140750 $D=0
M1367 184 1 4 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=145380 $D=0
M1368 2 173 182 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=136120 $D=0
M1369 3 174 183 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=140750 $D=0
M1370 4 175 184 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=145380 $D=0
M1371 188 5 182 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=136120 $D=0
M1372 189 5 183 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=140750 $D=0
M1373 190 5 184 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=145380 $D=0
M1374 185 5 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=136120 $D=0
M1375 186 5 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=140750 $D=0
M1376 187 5 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=145380 $D=0
M1377 191 5 179 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=136120 $D=0
M1378 192 5 180 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=140750 $D=0
M1379 193 5 181 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=145380 $D=0
M1380 176 185 191 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=136120 $D=0
M1381 177 186 192 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=140750 $D=0
M1382 178 187 193 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=145380 $D=0
M1383 194 6 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=136120 $D=0
M1384 195 6 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=140750 $D=0
M1385 196 6 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=145380 $D=0
M1386 197 6 191 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=136120 $D=0
M1387 198 6 192 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=140750 $D=0
M1388 199 6 193 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=145380 $D=0
M1389 188 194 197 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=136120 $D=0
M1390 189 195 198 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=140750 $D=0
M1391 190 196 199 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=145380 $D=0
M1392 200 7 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=136120 $D=0
M1393 201 7 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=140750 $D=0
M1394 202 7 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=145380 $D=0
M1395 203 7 8 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=136120 $D=0
M1396 204 7 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=140750 $D=0
M1397 205 7 10 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=145380 $D=0
M1398 11 200 203 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=136120 $D=0
M1399 12 201 204 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=140750 $D=0
M1400 13 202 205 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=145380 $D=0
M1401 206 7 14 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=136120 $D=0
M1402 207 7 15 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=140750 $D=0
M1403 208 7 16 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=145380 $D=0
M1404 209 200 206 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=136120 $D=0
M1405 210 201 207 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=140750 $D=0
M1406 211 202 208 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=145380 $D=0
M1407 215 7 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=136120 $D=0
M1408 216 7 213 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=140750 $D=0
M1409 217 7 214 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=145380 $D=0
M1410 197 200 215 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=136120 $D=0
M1411 198 201 216 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=140750 $D=0
M1412 199 202 217 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=145380 $D=0
M1413 221 17 215 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=136120 $D=0
M1414 222 17 216 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=140750 $D=0
M1415 223 17 217 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=145380 $D=0
M1416 218 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=136120 $D=0
M1417 219 17 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=140750 $D=0
M1418 220 17 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=145380 $D=0
M1419 224 17 206 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=136120 $D=0
M1420 225 17 207 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=140750 $D=0
M1421 226 17 208 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=145380 $D=0
M1422 203 218 224 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=136120 $D=0
M1423 204 219 225 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=140750 $D=0
M1424 205 220 226 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=145380 $D=0
M1425 227 18 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=136120 $D=0
M1426 228 18 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=140750 $D=0
M1427 229 18 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=145380 $D=0
M1428 230 18 224 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=136120 $D=0
M1429 231 18 225 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=140750 $D=0
M1430 232 18 226 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=145380 $D=0
M1431 221 227 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=136120 $D=0
M1432 222 228 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=140750 $D=0
M1433 223 229 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=145380 $D=0
M1434 167 19 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=136120 $D=0
M1435 171 19 234 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=140750 $D=0
M1436 172 19 235 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=145380 $D=0
M1437 236 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=136120 $D=0
M1438 237 20 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=140750 $D=0
M1439 238 20 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=145380 $D=0
M1440 239 233 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=136120 $D=0
M1441 240 234 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=140750 $D=0
M1442 241 235 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=145380 $D=0
M1443 167 239 940 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=136120 $D=0
M1444 171 240 941 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=140750 $D=0
M1445 172 241 942 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=145380 $D=0
M1446 242 940 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=136120 $D=0
M1447 243 941 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=140750 $D=0
M1448 244 942 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=145380 $D=0
M1449 239 19 242 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=136120 $D=0
M1450 240 19 243 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=140750 $D=0
M1451 241 19 244 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=145380 $D=0
M1452 242 236 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=136120 $D=0
M1453 243 237 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=140750 $D=0
M1454 244 238 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=145380 $D=0
M1455 251 248 242 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=136120 $D=0
M1456 252 249 243 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=140750 $D=0
M1457 253 250 244 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=145380 $D=0
M1458 248 21 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=136120 $D=0
M1459 249 21 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=140750 $D=0
M1460 250 21 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=145380 $D=0
M1461 167 22 254 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=136120 $D=0
M1462 171 22 255 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=140750 $D=0
M1463 172 22 256 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=145380 $D=0
M1464 257 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=136120 $D=0
M1465 258 23 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=140750 $D=0
M1466 259 23 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=145380 $D=0
M1467 260 254 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=136120 $D=0
M1468 261 255 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=140750 $D=0
M1469 262 256 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=145380 $D=0
M1470 167 260 943 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=136120 $D=0
M1471 171 261 944 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=140750 $D=0
M1472 172 262 945 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=145380 $D=0
M1473 263 943 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=136120 $D=0
M1474 264 944 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=140750 $D=0
M1475 265 945 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=145380 $D=0
M1476 260 22 263 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=136120 $D=0
M1477 261 22 264 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=140750 $D=0
M1478 262 22 265 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=145380 $D=0
M1479 263 257 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=136120 $D=0
M1480 264 258 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=140750 $D=0
M1481 265 259 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=145380 $D=0
M1482 251 266 263 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=136120 $D=0
M1483 252 267 264 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=140750 $D=0
M1484 253 268 265 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=145380 $D=0
M1485 266 24 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=136120 $D=0
M1486 267 24 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=140750 $D=0
M1487 268 24 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=145380 $D=0
M1488 167 25 269 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=136120 $D=0
M1489 171 25 270 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=140750 $D=0
M1490 172 25 271 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=145380 $D=0
M1491 272 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=136120 $D=0
M1492 273 26 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=140750 $D=0
M1493 274 26 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=145380 $D=0
M1494 275 269 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=136120 $D=0
M1495 276 270 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=140750 $D=0
M1496 277 271 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=145380 $D=0
M1497 167 275 946 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=136120 $D=0
M1498 171 276 947 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=140750 $D=0
M1499 172 277 948 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=145380 $D=0
M1500 278 946 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=136120 $D=0
M1501 279 947 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=140750 $D=0
M1502 280 948 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=145380 $D=0
M1503 275 25 278 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=136120 $D=0
M1504 276 25 279 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=140750 $D=0
M1505 277 25 280 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=145380 $D=0
M1506 278 272 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=136120 $D=0
M1507 279 273 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=140750 $D=0
M1508 280 274 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=145380 $D=0
M1509 251 281 278 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=136120 $D=0
M1510 252 282 279 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=140750 $D=0
M1511 253 283 280 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=145380 $D=0
M1512 281 27 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=136120 $D=0
M1513 282 27 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=140750 $D=0
M1514 283 27 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=145380 $D=0
M1515 167 28 284 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=136120 $D=0
M1516 171 28 285 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=140750 $D=0
M1517 172 28 286 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=145380 $D=0
M1518 287 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=136120 $D=0
M1519 288 29 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=140750 $D=0
M1520 289 29 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=145380 $D=0
M1521 290 284 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=136120 $D=0
M1522 291 285 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=140750 $D=0
M1523 292 286 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=145380 $D=0
M1524 167 290 949 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=136120 $D=0
M1525 171 291 950 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=140750 $D=0
M1526 172 292 951 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=145380 $D=0
M1527 293 949 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=136120 $D=0
M1528 294 950 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=140750 $D=0
M1529 295 951 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=145380 $D=0
M1530 290 28 293 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=136120 $D=0
M1531 291 28 294 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=140750 $D=0
M1532 292 28 295 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=145380 $D=0
M1533 293 287 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=136120 $D=0
M1534 294 288 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=140750 $D=0
M1535 295 289 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=145380 $D=0
M1536 251 296 293 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=136120 $D=0
M1537 252 297 294 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=140750 $D=0
M1538 253 298 295 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=145380 $D=0
M1539 296 30 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=136120 $D=0
M1540 297 30 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=140750 $D=0
M1541 298 30 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=145380 $D=0
M1542 167 31 299 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=136120 $D=0
M1543 171 31 300 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=140750 $D=0
M1544 172 31 301 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=145380 $D=0
M1545 302 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=136120 $D=0
M1546 303 32 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=140750 $D=0
M1547 304 32 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=145380 $D=0
M1548 305 299 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=136120 $D=0
M1549 306 300 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=140750 $D=0
M1550 307 301 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=145380 $D=0
M1551 167 305 952 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=136120 $D=0
M1552 171 306 953 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=140750 $D=0
M1553 172 307 954 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=145380 $D=0
M1554 308 952 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=136120 $D=0
M1555 309 953 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=140750 $D=0
M1556 310 954 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=145380 $D=0
M1557 305 31 308 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=136120 $D=0
M1558 306 31 309 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=140750 $D=0
M1559 307 31 310 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=145380 $D=0
M1560 308 302 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=136120 $D=0
M1561 309 303 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=140750 $D=0
M1562 310 304 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=145380 $D=0
M1563 251 311 308 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=136120 $D=0
M1564 252 312 309 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=140750 $D=0
M1565 253 313 310 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=145380 $D=0
M1566 311 33 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=136120 $D=0
M1567 312 33 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=140750 $D=0
M1568 313 33 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=145380 $D=0
M1569 167 34 314 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=136120 $D=0
M1570 171 34 315 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=140750 $D=0
M1571 172 34 316 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=145380 $D=0
M1572 317 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=136120 $D=0
M1573 318 35 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=140750 $D=0
M1574 319 35 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=145380 $D=0
M1575 320 314 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=136120 $D=0
M1576 321 315 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=140750 $D=0
M1577 322 316 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=145380 $D=0
M1578 167 320 955 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=136120 $D=0
M1579 171 321 956 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=140750 $D=0
M1580 172 322 957 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=145380 $D=0
M1581 323 955 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=136120 $D=0
M1582 324 956 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=140750 $D=0
M1583 325 957 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=145380 $D=0
M1584 320 34 323 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=136120 $D=0
M1585 321 34 324 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=140750 $D=0
M1586 322 34 325 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=145380 $D=0
M1587 323 317 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=136120 $D=0
M1588 324 318 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=140750 $D=0
M1589 325 319 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=145380 $D=0
M1590 251 326 323 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=136120 $D=0
M1591 252 327 324 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=140750 $D=0
M1592 253 328 325 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=145380 $D=0
M1593 326 36 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=136120 $D=0
M1594 327 36 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=140750 $D=0
M1595 328 36 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=145380 $D=0
M1596 167 37 329 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=136120 $D=0
M1597 171 37 330 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=140750 $D=0
M1598 172 37 331 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=145380 $D=0
M1599 332 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=136120 $D=0
M1600 333 38 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=140750 $D=0
M1601 334 38 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=145380 $D=0
M1602 335 329 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=136120 $D=0
M1603 336 330 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=140750 $D=0
M1604 337 331 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=145380 $D=0
M1605 167 335 958 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=136120 $D=0
M1606 171 336 959 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=140750 $D=0
M1607 172 337 960 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=145380 $D=0
M1608 338 958 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=136120 $D=0
M1609 339 959 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=140750 $D=0
M1610 340 960 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=145380 $D=0
M1611 335 37 338 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=136120 $D=0
M1612 336 37 339 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=140750 $D=0
M1613 337 37 340 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=145380 $D=0
M1614 338 332 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=136120 $D=0
M1615 339 333 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=140750 $D=0
M1616 340 334 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=145380 $D=0
M1617 251 341 338 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=136120 $D=0
M1618 252 342 339 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=140750 $D=0
M1619 253 343 340 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=145380 $D=0
M1620 341 39 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=136120 $D=0
M1621 342 39 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=140750 $D=0
M1622 343 39 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=145380 $D=0
M1623 167 40 344 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=136120 $D=0
M1624 171 40 345 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=140750 $D=0
M1625 172 40 346 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=145380 $D=0
M1626 347 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=136120 $D=0
M1627 348 41 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=140750 $D=0
M1628 349 41 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=145380 $D=0
M1629 350 344 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=136120 $D=0
M1630 351 345 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=140750 $D=0
M1631 352 346 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=145380 $D=0
M1632 167 350 961 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=136120 $D=0
M1633 171 351 962 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=140750 $D=0
M1634 172 352 963 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=145380 $D=0
M1635 353 961 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=136120 $D=0
M1636 354 962 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=140750 $D=0
M1637 355 963 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=145380 $D=0
M1638 350 40 353 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=136120 $D=0
M1639 351 40 354 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=140750 $D=0
M1640 352 40 355 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=145380 $D=0
M1641 353 347 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=136120 $D=0
M1642 354 348 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=140750 $D=0
M1643 355 349 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=145380 $D=0
M1644 251 356 353 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=136120 $D=0
M1645 252 357 354 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=140750 $D=0
M1646 253 358 355 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=145380 $D=0
M1647 356 42 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=136120 $D=0
M1648 357 42 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=140750 $D=0
M1649 358 42 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=145380 $D=0
M1650 167 43 359 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=136120 $D=0
M1651 171 43 360 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=140750 $D=0
M1652 172 43 361 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=145380 $D=0
M1653 362 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=136120 $D=0
M1654 363 44 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=140750 $D=0
M1655 364 44 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=145380 $D=0
M1656 365 359 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=136120 $D=0
M1657 366 360 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=140750 $D=0
M1658 367 361 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=145380 $D=0
M1659 167 365 964 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=136120 $D=0
M1660 171 366 965 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=140750 $D=0
M1661 172 367 966 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=145380 $D=0
M1662 368 964 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=136120 $D=0
M1663 369 965 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=140750 $D=0
M1664 370 966 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=145380 $D=0
M1665 365 43 368 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=136120 $D=0
M1666 366 43 369 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=140750 $D=0
M1667 367 43 370 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=145380 $D=0
M1668 368 362 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=136120 $D=0
M1669 369 363 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=140750 $D=0
M1670 370 364 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=145380 $D=0
M1671 251 371 368 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=136120 $D=0
M1672 252 372 369 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=140750 $D=0
M1673 253 373 370 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=145380 $D=0
M1674 371 45 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=136120 $D=0
M1675 372 45 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=140750 $D=0
M1676 373 45 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=145380 $D=0
M1677 167 46 374 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=136120 $D=0
M1678 171 46 375 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=140750 $D=0
M1679 172 46 376 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=145380 $D=0
M1680 377 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=136120 $D=0
M1681 378 47 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=140750 $D=0
M1682 379 47 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=145380 $D=0
M1683 380 374 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=136120 $D=0
M1684 381 375 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=140750 $D=0
M1685 382 376 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=145380 $D=0
M1686 167 380 967 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=136120 $D=0
M1687 171 381 968 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=140750 $D=0
M1688 172 382 969 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=145380 $D=0
M1689 383 967 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=136120 $D=0
M1690 384 968 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=140750 $D=0
M1691 385 969 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=145380 $D=0
M1692 380 46 383 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=136120 $D=0
M1693 381 46 384 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=140750 $D=0
M1694 382 46 385 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=145380 $D=0
M1695 383 377 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=136120 $D=0
M1696 384 378 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=140750 $D=0
M1697 385 379 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=145380 $D=0
M1698 251 386 383 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=136120 $D=0
M1699 252 387 384 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=140750 $D=0
M1700 253 388 385 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=145380 $D=0
M1701 386 48 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=136120 $D=0
M1702 387 48 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=140750 $D=0
M1703 388 48 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=145380 $D=0
M1704 167 49 389 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=136120 $D=0
M1705 171 49 390 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=140750 $D=0
M1706 172 49 391 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=145380 $D=0
M1707 392 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=136120 $D=0
M1708 393 50 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=140750 $D=0
M1709 394 50 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=145380 $D=0
M1710 395 389 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=136120 $D=0
M1711 396 390 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=140750 $D=0
M1712 397 391 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=145380 $D=0
M1713 167 395 970 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=136120 $D=0
M1714 171 396 971 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=140750 $D=0
M1715 172 397 972 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=145380 $D=0
M1716 398 970 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=136120 $D=0
M1717 399 971 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=140750 $D=0
M1718 400 972 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=145380 $D=0
M1719 395 49 398 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=136120 $D=0
M1720 396 49 399 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=140750 $D=0
M1721 397 49 400 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=145380 $D=0
M1722 398 392 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=136120 $D=0
M1723 399 393 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=140750 $D=0
M1724 400 394 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=145380 $D=0
M1725 251 401 398 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=136120 $D=0
M1726 252 402 399 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=140750 $D=0
M1727 253 403 400 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=145380 $D=0
M1728 401 51 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=136120 $D=0
M1729 402 51 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=140750 $D=0
M1730 403 51 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=145380 $D=0
M1731 167 52 404 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=136120 $D=0
M1732 171 52 405 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=140750 $D=0
M1733 172 52 406 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=145380 $D=0
M1734 407 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=136120 $D=0
M1735 408 53 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=140750 $D=0
M1736 409 53 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=145380 $D=0
M1737 410 404 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=136120 $D=0
M1738 411 405 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=140750 $D=0
M1739 412 406 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=145380 $D=0
M1740 167 410 973 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=136120 $D=0
M1741 171 411 974 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=140750 $D=0
M1742 172 412 975 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=145380 $D=0
M1743 413 973 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=136120 $D=0
M1744 414 974 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=140750 $D=0
M1745 415 975 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=145380 $D=0
M1746 410 52 413 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=136120 $D=0
M1747 411 52 414 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=140750 $D=0
M1748 412 52 415 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=145380 $D=0
M1749 413 407 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=136120 $D=0
M1750 414 408 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=140750 $D=0
M1751 415 409 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=145380 $D=0
M1752 251 416 413 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=136120 $D=0
M1753 252 417 414 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=140750 $D=0
M1754 253 418 415 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=145380 $D=0
M1755 416 54 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=136120 $D=0
M1756 417 54 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=140750 $D=0
M1757 418 54 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=145380 $D=0
M1758 167 55 419 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=136120 $D=0
M1759 171 55 420 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=140750 $D=0
M1760 172 55 421 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=145380 $D=0
M1761 422 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=136120 $D=0
M1762 423 56 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=140750 $D=0
M1763 424 56 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=145380 $D=0
M1764 425 419 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=136120 $D=0
M1765 426 420 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=140750 $D=0
M1766 427 421 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=145380 $D=0
M1767 167 425 976 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=136120 $D=0
M1768 171 426 977 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=140750 $D=0
M1769 172 427 978 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=145380 $D=0
M1770 428 976 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=136120 $D=0
M1771 429 977 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=140750 $D=0
M1772 430 978 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=145380 $D=0
M1773 425 55 428 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=136120 $D=0
M1774 426 55 429 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=140750 $D=0
M1775 427 55 430 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=145380 $D=0
M1776 428 422 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=136120 $D=0
M1777 429 423 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=140750 $D=0
M1778 430 424 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=145380 $D=0
M1779 251 431 428 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=136120 $D=0
M1780 252 432 429 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=140750 $D=0
M1781 253 433 430 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=145380 $D=0
M1782 431 57 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=136120 $D=0
M1783 432 57 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=140750 $D=0
M1784 433 57 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=145380 $D=0
M1785 167 58 434 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=136120 $D=0
M1786 171 58 435 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=140750 $D=0
M1787 172 58 436 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=145380 $D=0
M1788 437 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=136120 $D=0
M1789 438 59 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=140750 $D=0
M1790 439 59 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=145380 $D=0
M1791 440 434 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=136120 $D=0
M1792 441 435 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=140750 $D=0
M1793 442 436 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=145380 $D=0
M1794 167 440 979 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=136120 $D=0
M1795 171 441 980 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=140750 $D=0
M1796 172 442 981 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=145380 $D=0
M1797 443 979 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=136120 $D=0
M1798 444 980 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=140750 $D=0
M1799 445 981 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=145380 $D=0
M1800 440 58 443 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=136120 $D=0
M1801 441 58 444 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=140750 $D=0
M1802 442 58 445 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=145380 $D=0
M1803 443 437 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=136120 $D=0
M1804 444 438 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=140750 $D=0
M1805 445 439 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=145380 $D=0
M1806 251 446 443 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=136120 $D=0
M1807 252 447 444 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=140750 $D=0
M1808 253 448 445 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=145380 $D=0
M1809 446 60 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=136120 $D=0
M1810 447 60 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=140750 $D=0
M1811 448 60 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=145380 $D=0
M1812 167 61 449 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=136120 $D=0
M1813 171 61 450 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=140750 $D=0
M1814 172 61 451 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=145380 $D=0
M1815 452 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=136120 $D=0
M1816 453 62 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=140750 $D=0
M1817 454 62 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=145380 $D=0
M1818 455 449 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=136120 $D=0
M1819 456 450 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=140750 $D=0
M1820 457 451 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=145380 $D=0
M1821 167 455 982 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=136120 $D=0
M1822 171 456 983 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=140750 $D=0
M1823 172 457 984 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=145380 $D=0
M1824 458 982 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=136120 $D=0
M1825 459 983 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=140750 $D=0
M1826 460 984 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=145380 $D=0
M1827 455 61 458 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=136120 $D=0
M1828 456 61 459 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=140750 $D=0
M1829 457 61 460 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=145380 $D=0
M1830 458 452 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=136120 $D=0
M1831 459 453 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=140750 $D=0
M1832 460 454 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=145380 $D=0
M1833 251 461 458 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=136120 $D=0
M1834 252 462 459 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=140750 $D=0
M1835 253 463 460 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=145380 $D=0
M1836 461 63 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=136120 $D=0
M1837 462 63 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=140750 $D=0
M1838 463 63 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=145380 $D=0
M1839 167 64 464 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=136120 $D=0
M1840 171 64 465 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=140750 $D=0
M1841 172 64 466 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=145380 $D=0
M1842 467 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=136120 $D=0
M1843 468 65 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=140750 $D=0
M1844 469 65 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=145380 $D=0
M1845 470 464 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=136120 $D=0
M1846 471 465 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=140750 $D=0
M1847 472 466 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=145380 $D=0
M1848 167 470 985 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=136120 $D=0
M1849 171 471 986 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=140750 $D=0
M1850 172 472 987 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=145380 $D=0
M1851 473 985 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=136120 $D=0
M1852 474 986 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=140750 $D=0
M1853 475 987 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=145380 $D=0
M1854 470 64 473 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=136120 $D=0
M1855 471 64 474 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=140750 $D=0
M1856 472 64 475 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=145380 $D=0
M1857 473 467 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=136120 $D=0
M1858 474 468 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=140750 $D=0
M1859 475 469 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=145380 $D=0
M1860 251 476 473 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=136120 $D=0
M1861 252 477 474 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=140750 $D=0
M1862 253 478 475 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=145380 $D=0
M1863 476 66 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=136120 $D=0
M1864 477 66 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=140750 $D=0
M1865 478 66 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=145380 $D=0
M1866 167 67 479 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=136120 $D=0
M1867 171 67 480 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=140750 $D=0
M1868 172 67 481 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=145380 $D=0
M1869 482 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=136120 $D=0
M1870 483 68 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=140750 $D=0
M1871 484 68 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=145380 $D=0
M1872 485 479 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=136120 $D=0
M1873 486 480 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=140750 $D=0
M1874 487 481 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=145380 $D=0
M1875 167 485 988 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=136120 $D=0
M1876 171 486 989 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=140750 $D=0
M1877 172 487 990 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=145380 $D=0
M1878 488 988 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=136120 $D=0
M1879 489 989 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=140750 $D=0
M1880 490 990 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=145380 $D=0
M1881 485 67 488 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=136120 $D=0
M1882 486 67 489 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=140750 $D=0
M1883 487 67 490 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=145380 $D=0
M1884 488 482 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=136120 $D=0
M1885 489 483 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=140750 $D=0
M1886 490 484 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=145380 $D=0
M1887 251 491 488 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=136120 $D=0
M1888 252 492 489 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=140750 $D=0
M1889 253 493 490 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=145380 $D=0
M1890 491 69 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=136120 $D=0
M1891 492 69 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=140750 $D=0
M1892 493 69 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=145380 $D=0
M1893 167 70 494 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=136120 $D=0
M1894 171 70 495 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=140750 $D=0
M1895 172 70 496 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=145380 $D=0
M1896 497 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=136120 $D=0
M1897 498 71 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=140750 $D=0
M1898 499 71 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=145380 $D=0
M1899 500 494 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=136120 $D=0
M1900 501 495 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=140750 $D=0
M1901 502 496 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=145380 $D=0
M1902 167 500 991 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=136120 $D=0
M1903 171 501 992 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=140750 $D=0
M1904 172 502 993 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=145380 $D=0
M1905 503 991 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=136120 $D=0
M1906 504 992 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=140750 $D=0
M1907 505 993 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=145380 $D=0
M1908 500 70 503 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=136120 $D=0
M1909 501 70 504 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=140750 $D=0
M1910 502 70 505 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=145380 $D=0
M1911 503 497 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=136120 $D=0
M1912 504 498 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=140750 $D=0
M1913 505 499 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=145380 $D=0
M1914 251 506 503 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=136120 $D=0
M1915 252 507 504 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=140750 $D=0
M1916 253 508 505 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=145380 $D=0
M1917 506 72 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=136120 $D=0
M1918 507 72 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=140750 $D=0
M1919 508 72 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=145380 $D=0
M1920 167 73 509 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=136120 $D=0
M1921 171 73 510 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=140750 $D=0
M1922 172 73 511 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=145380 $D=0
M1923 512 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=136120 $D=0
M1924 513 74 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=140750 $D=0
M1925 514 74 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=145380 $D=0
M1926 515 509 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=136120 $D=0
M1927 516 510 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=140750 $D=0
M1928 517 511 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=145380 $D=0
M1929 167 515 994 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=136120 $D=0
M1930 171 516 995 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=140750 $D=0
M1931 172 517 996 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=145380 $D=0
M1932 518 994 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=136120 $D=0
M1933 519 995 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=140750 $D=0
M1934 520 996 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=145380 $D=0
M1935 515 73 518 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=136120 $D=0
M1936 516 73 519 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=140750 $D=0
M1937 517 73 520 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=145380 $D=0
M1938 518 512 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=136120 $D=0
M1939 519 513 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=140750 $D=0
M1940 520 514 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=145380 $D=0
M1941 251 521 518 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=136120 $D=0
M1942 252 522 519 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=140750 $D=0
M1943 253 523 520 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=145380 $D=0
M1944 521 75 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=136120 $D=0
M1945 522 75 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=140750 $D=0
M1946 523 75 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=145380 $D=0
M1947 167 76 524 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=136120 $D=0
M1948 171 76 525 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=140750 $D=0
M1949 172 76 526 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=145380 $D=0
M1950 527 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=136120 $D=0
M1951 528 77 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=140750 $D=0
M1952 529 77 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=145380 $D=0
M1953 530 524 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=136120 $D=0
M1954 531 525 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=140750 $D=0
M1955 532 526 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=145380 $D=0
M1956 167 530 997 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=136120 $D=0
M1957 171 531 998 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=140750 $D=0
M1958 172 532 999 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=145380 $D=0
M1959 533 997 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=136120 $D=0
M1960 534 998 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=140750 $D=0
M1961 535 999 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=145380 $D=0
M1962 530 76 533 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=136120 $D=0
M1963 531 76 534 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=140750 $D=0
M1964 532 76 535 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=145380 $D=0
M1965 533 527 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=136120 $D=0
M1966 534 528 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=140750 $D=0
M1967 535 529 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=145380 $D=0
M1968 251 536 533 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=136120 $D=0
M1969 252 537 534 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=140750 $D=0
M1970 253 538 535 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=145380 $D=0
M1971 536 78 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=136120 $D=0
M1972 537 78 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=140750 $D=0
M1973 538 78 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=145380 $D=0
M1974 167 79 539 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=136120 $D=0
M1975 171 79 540 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=140750 $D=0
M1976 172 79 541 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=145380 $D=0
M1977 542 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=136120 $D=0
M1978 543 80 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=140750 $D=0
M1979 544 80 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=145380 $D=0
M1980 545 539 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=136120 $D=0
M1981 546 540 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=140750 $D=0
M1982 547 541 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=145380 $D=0
M1983 167 545 1000 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=136120 $D=0
M1984 171 546 1001 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=140750 $D=0
M1985 172 547 1002 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=145380 $D=0
M1986 548 1000 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=136120 $D=0
M1987 549 1001 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=140750 $D=0
M1988 550 1002 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=145380 $D=0
M1989 545 79 548 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=136120 $D=0
M1990 546 79 549 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=140750 $D=0
M1991 547 79 550 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=145380 $D=0
M1992 548 542 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=136120 $D=0
M1993 549 543 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=140750 $D=0
M1994 550 544 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=145380 $D=0
M1995 251 551 548 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=136120 $D=0
M1996 252 552 549 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=140750 $D=0
M1997 253 553 550 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=145380 $D=0
M1998 551 81 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=136120 $D=0
M1999 552 81 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=140750 $D=0
M2000 553 81 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=145380 $D=0
M2001 167 82 554 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=136120 $D=0
M2002 171 82 555 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=140750 $D=0
M2003 172 82 556 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=145380 $D=0
M2004 557 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=136120 $D=0
M2005 558 83 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=140750 $D=0
M2006 559 83 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=145380 $D=0
M2007 560 554 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=136120 $D=0
M2008 561 555 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=140750 $D=0
M2009 562 556 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=145380 $D=0
M2010 167 560 1003 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=136120 $D=0
M2011 171 561 1004 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=140750 $D=0
M2012 172 562 1005 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=145380 $D=0
M2013 563 1003 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=136120 $D=0
M2014 564 1004 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=140750 $D=0
M2015 565 1005 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=145380 $D=0
M2016 560 82 563 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=136120 $D=0
M2017 561 82 564 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=140750 $D=0
M2018 562 82 565 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=145380 $D=0
M2019 563 557 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=136120 $D=0
M2020 564 558 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=140750 $D=0
M2021 565 559 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=145380 $D=0
M2022 251 566 563 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=136120 $D=0
M2023 252 567 564 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=140750 $D=0
M2024 253 568 565 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=145380 $D=0
M2025 566 84 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=136120 $D=0
M2026 567 84 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=140750 $D=0
M2027 568 84 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=145380 $D=0
M2028 167 85 569 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=136120 $D=0
M2029 171 85 570 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=140750 $D=0
M2030 172 85 571 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=145380 $D=0
M2031 572 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=136120 $D=0
M2032 573 86 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=140750 $D=0
M2033 574 86 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=145380 $D=0
M2034 575 569 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=136120 $D=0
M2035 576 570 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=140750 $D=0
M2036 577 571 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=145380 $D=0
M2037 167 575 1006 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=136120 $D=0
M2038 171 576 1007 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=140750 $D=0
M2039 172 577 1008 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=145380 $D=0
M2040 578 1006 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=136120 $D=0
M2041 579 1007 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=140750 $D=0
M2042 580 1008 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=145380 $D=0
M2043 575 85 578 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=136120 $D=0
M2044 576 85 579 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=140750 $D=0
M2045 577 85 580 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=145380 $D=0
M2046 578 572 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=136120 $D=0
M2047 579 573 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=140750 $D=0
M2048 580 574 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=145380 $D=0
M2049 251 581 578 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=136120 $D=0
M2050 252 582 579 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=140750 $D=0
M2051 253 583 580 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=145380 $D=0
M2052 581 87 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=136120 $D=0
M2053 582 87 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=140750 $D=0
M2054 583 87 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=145380 $D=0
M2055 167 88 584 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=136120 $D=0
M2056 171 88 585 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=140750 $D=0
M2057 172 88 586 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=145380 $D=0
M2058 587 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=136120 $D=0
M2059 588 89 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=140750 $D=0
M2060 589 89 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=145380 $D=0
M2061 590 584 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=136120 $D=0
M2062 591 585 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=140750 $D=0
M2063 592 586 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=145380 $D=0
M2064 167 590 1009 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=136120 $D=0
M2065 171 591 1010 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=140750 $D=0
M2066 172 592 1011 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=145380 $D=0
M2067 593 1009 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=136120 $D=0
M2068 594 1010 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=140750 $D=0
M2069 595 1011 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=145380 $D=0
M2070 590 88 593 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=136120 $D=0
M2071 591 88 594 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=140750 $D=0
M2072 592 88 595 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=145380 $D=0
M2073 593 587 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=136120 $D=0
M2074 594 588 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=140750 $D=0
M2075 595 589 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=145380 $D=0
M2076 251 596 593 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=136120 $D=0
M2077 252 597 594 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=140750 $D=0
M2078 253 598 595 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=145380 $D=0
M2079 596 90 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=136120 $D=0
M2080 597 90 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=140750 $D=0
M2081 598 90 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=145380 $D=0
M2082 167 91 599 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=136120 $D=0
M2083 171 91 600 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=140750 $D=0
M2084 172 91 601 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=145380 $D=0
M2085 602 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=136120 $D=0
M2086 603 92 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=140750 $D=0
M2087 604 92 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=145380 $D=0
M2088 605 599 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=136120 $D=0
M2089 606 600 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=140750 $D=0
M2090 607 601 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=145380 $D=0
M2091 167 605 1012 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=136120 $D=0
M2092 171 606 1013 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=140750 $D=0
M2093 172 607 1014 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=145380 $D=0
M2094 608 1012 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=136120 $D=0
M2095 609 1013 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=140750 $D=0
M2096 610 1014 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=145380 $D=0
M2097 605 91 608 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=136120 $D=0
M2098 606 91 609 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=140750 $D=0
M2099 607 91 610 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=145380 $D=0
M2100 608 602 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=136120 $D=0
M2101 609 603 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=140750 $D=0
M2102 610 604 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=145380 $D=0
M2103 251 611 608 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=136120 $D=0
M2104 252 612 609 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=140750 $D=0
M2105 253 613 610 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=145380 $D=0
M2106 611 93 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=136120 $D=0
M2107 612 93 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=140750 $D=0
M2108 613 93 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=145380 $D=0
M2109 167 94 614 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=136120 $D=0
M2110 171 94 615 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=140750 $D=0
M2111 172 94 616 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=145380 $D=0
M2112 617 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=136120 $D=0
M2113 618 95 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=140750 $D=0
M2114 619 95 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=145380 $D=0
M2115 620 614 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=136120 $D=0
M2116 621 615 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=140750 $D=0
M2117 622 616 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=145380 $D=0
M2118 167 620 1015 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=136120 $D=0
M2119 171 621 1016 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=140750 $D=0
M2120 172 622 1017 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=145380 $D=0
M2121 623 1015 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=136120 $D=0
M2122 624 1016 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=140750 $D=0
M2123 625 1017 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=145380 $D=0
M2124 620 94 623 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=136120 $D=0
M2125 621 94 624 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=140750 $D=0
M2126 622 94 625 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=145380 $D=0
M2127 623 617 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=136120 $D=0
M2128 624 618 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=140750 $D=0
M2129 625 619 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=145380 $D=0
M2130 251 626 623 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=136120 $D=0
M2131 252 627 624 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=140750 $D=0
M2132 253 628 625 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=145380 $D=0
M2133 626 96 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=136120 $D=0
M2134 627 96 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=140750 $D=0
M2135 628 96 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=145380 $D=0
M2136 167 97 629 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=136120 $D=0
M2137 171 97 630 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=140750 $D=0
M2138 172 97 631 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=145380 $D=0
M2139 632 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=136120 $D=0
M2140 633 98 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=140750 $D=0
M2141 634 98 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=145380 $D=0
M2142 635 629 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=136120 $D=0
M2143 636 630 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=140750 $D=0
M2144 637 631 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=145380 $D=0
M2145 167 635 1018 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=136120 $D=0
M2146 171 636 1019 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=140750 $D=0
M2147 172 637 1020 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=145380 $D=0
M2148 638 1018 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=136120 $D=0
M2149 639 1019 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=140750 $D=0
M2150 640 1020 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=145380 $D=0
M2151 635 97 638 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=136120 $D=0
M2152 636 97 639 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=140750 $D=0
M2153 637 97 640 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=145380 $D=0
M2154 638 632 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=136120 $D=0
M2155 639 633 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=140750 $D=0
M2156 640 634 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=145380 $D=0
M2157 251 641 638 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=136120 $D=0
M2158 252 642 639 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=140750 $D=0
M2159 253 643 640 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=145380 $D=0
M2160 641 99 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=136120 $D=0
M2161 642 99 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=140750 $D=0
M2162 643 99 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=145380 $D=0
M2163 167 100 644 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=136120 $D=0
M2164 171 100 645 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=140750 $D=0
M2165 172 100 646 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=145380 $D=0
M2166 647 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=136120 $D=0
M2167 648 101 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=140750 $D=0
M2168 649 101 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=145380 $D=0
M2169 650 644 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=136120 $D=0
M2170 651 645 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=140750 $D=0
M2171 652 646 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=145380 $D=0
M2172 167 650 1021 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=136120 $D=0
M2173 171 651 1022 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=140750 $D=0
M2174 172 652 1023 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=145380 $D=0
M2175 653 1021 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=136120 $D=0
M2176 654 1022 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=140750 $D=0
M2177 655 1023 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=145380 $D=0
M2178 650 100 653 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=136120 $D=0
M2179 651 100 654 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=140750 $D=0
M2180 652 100 655 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=145380 $D=0
M2181 653 647 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=136120 $D=0
M2182 654 648 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=140750 $D=0
M2183 655 649 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=145380 $D=0
M2184 251 656 653 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=136120 $D=0
M2185 252 657 654 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=140750 $D=0
M2186 253 658 655 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=145380 $D=0
M2187 656 102 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=136120 $D=0
M2188 657 102 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=140750 $D=0
M2189 658 102 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=145380 $D=0
M2190 167 103 659 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=136120 $D=0
M2191 171 103 660 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=140750 $D=0
M2192 172 103 661 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=145380 $D=0
M2193 662 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=136120 $D=0
M2194 663 104 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=140750 $D=0
M2195 664 104 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=145380 $D=0
M2196 665 659 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=136120 $D=0
M2197 666 660 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=140750 $D=0
M2198 667 661 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=145380 $D=0
M2199 167 665 1024 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=136120 $D=0
M2200 171 666 1025 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=140750 $D=0
M2201 172 667 1026 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=145380 $D=0
M2202 668 1024 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=136120 $D=0
M2203 669 1025 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=140750 $D=0
M2204 670 1026 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=145380 $D=0
M2205 665 103 668 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=136120 $D=0
M2206 666 103 669 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=140750 $D=0
M2207 667 103 670 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=145380 $D=0
M2208 668 662 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=136120 $D=0
M2209 669 663 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=140750 $D=0
M2210 670 664 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=145380 $D=0
M2211 251 671 668 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=136120 $D=0
M2212 252 672 669 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=140750 $D=0
M2213 253 673 670 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=145380 $D=0
M2214 671 105 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=136120 $D=0
M2215 672 105 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=140750 $D=0
M2216 673 105 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=145380 $D=0
M2217 167 106 674 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=136120 $D=0
M2218 171 106 675 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=140750 $D=0
M2219 172 106 676 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=145380 $D=0
M2220 677 107 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=136120 $D=0
M2221 678 107 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=140750 $D=0
M2222 679 107 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=145380 $D=0
M2223 680 674 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=136120 $D=0
M2224 681 675 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=140750 $D=0
M2225 682 676 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=145380 $D=0
M2226 167 680 1027 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=136120 $D=0
M2227 171 681 1028 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=140750 $D=0
M2228 172 682 1029 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=145380 $D=0
M2229 683 1027 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=136120 $D=0
M2230 684 1028 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=140750 $D=0
M2231 685 1029 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=145380 $D=0
M2232 680 106 683 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=136120 $D=0
M2233 681 106 684 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=140750 $D=0
M2234 682 106 685 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=145380 $D=0
M2235 683 677 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=136120 $D=0
M2236 684 678 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=140750 $D=0
M2237 685 679 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=145380 $D=0
M2238 251 686 683 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=136120 $D=0
M2239 252 687 684 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=140750 $D=0
M2240 253 688 685 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=145380 $D=0
M2241 686 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=136120 $D=0
M2242 687 108 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=140750 $D=0
M2243 688 108 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=145380 $D=0
M2244 167 109 689 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=136120 $D=0
M2245 171 109 690 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=140750 $D=0
M2246 172 109 691 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=145380 $D=0
M2247 692 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=136120 $D=0
M2248 693 110 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=140750 $D=0
M2249 694 110 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=145380 $D=0
M2250 695 689 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=136120 $D=0
M2251 696 690 231 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=140750 $D=0
M2252 697 691 232 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=145380 $D=0
M2253 167 695 1030 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=136120 $D=0
M2254 171 696 1031 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=140750 $D=0
M2255 172 697 1032 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=145380 $D=0
M2256 698 1030 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=136120 $D=0
M2257 699 1031 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=140750 $D=0
M2258 700 1032 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=145380 $D=0
M2259 695 109 698 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=136120 $D=0
M2260 696 109 699 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=140750 $D=0
M2261 697 109 700 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=145380 $D=0
M2262 698 692 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=136120 $D=0
M2263 699 693 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=140750 $D=0
M2264 700 694 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=145380 $D=0
M2265 251 701 698 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=136120 $D=0
M2266 252 702 699 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=140750 $D=0
M2267 253 703 700 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=145380 $D=0
M2268 701 111 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=136120 $D=0
M2269 702 111 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=140750 $D=0
M2270 703 111 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=145380 $D=0
M2271 167 112 704 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=136120 $D=0
M2272 171 112 705 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=140750 $D=0
M2273 172 112 706 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=145380 $D=0
M2274 707 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=136120 $D=0
M2275 708 113 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=140750 $D=0
M2276 709 113 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=145380 $D=0
M2277 8 707 245 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=136120 $D=0
M2278 9 708 246 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=140750 $D=0
M2279 140 709 247 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=145380 $D=0
M2280 251 704 8 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=136120 $D=0
M2281 252 705 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=140750 $D=0
M2282 253 706 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=145380 $D=0
M2283 167 713 710 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=136120 $D=0
M2284 171 714 711 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=140750 $D=0
M2285 172 715 712 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=145380 $D=0
M2286 713 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=136120 $D=0
M2287 714 114 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=140750 $D=0
M2288 715 114 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=145380 $D=0
M2289 1033 245 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=136120 $D=0
M2290 1034 246 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=140750 $D=0
M2291 1035 247 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=145380 $D=0
M2292 716 713 1033 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=136120 $D=0
M2293 717 714 1034 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=140750 $D=0
M2294 718 715 1035 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=145380 $D=0
M2295 167 716 719 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=136120 $D=0
M2296 171 717 720 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=140750 $D=0
M2297 172 718 721 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=145380 $D=0
M2298 1036 719 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=136120 $D=0
M2299 1037 720 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=140750 $D=0
M2300 1038 721 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=145380 $D=0
M2301 716 710 1036 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=136120 $D=0
M2302 717 711 1037 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=140750 $D=0
M2303 718 712 1038 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=145380 $D=0
M2304 167 725 722 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=136120 $D=0
M2305 171 726 723 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=140750 $D=0
M2306 172 727 724 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=145380 $D=0
M2307 725 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=136120 $D=0
M2308 726 114 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=140750 $D=0
M2309 727 114 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=145380 $D=0
M2310 1039 251 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=136120 $D=0
M2311 1040 252 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=140750 $D=0
M2312 1041 253 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=145380 $D=0
M2313 728 725 1039 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=136120 $D=0
M2314 729 726 1040 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=140750 $D=0
M2315 730 727 1041 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=145380 $D=0
M2316 167 728 115 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=136120 $D=0
M2317 171 729 116 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=140750 $D=0
M2318 172 730 117 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=145380 $D=0
M2319 1042 115 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=136120 $D=0
M2320 1043 116 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=140750 $D=0
M2321 1044 117 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=145380 $D=0
M2322 728 722 1042 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=136120 $D=0
M2323 729 723 1043 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=140750 $D=0
M2324 730 724 1044 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=145380 $D=0
M2325 731 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=136120 $D=0
M2326 732 118 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=140750 $D=0
M2327 733 118 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=145380 $D=0
M2328 734 118 719 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=136120 $D=0
M2329 735 118 720 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=140750 $D=0
M2330 736 118 721 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=145380 $D=0
M2331 119 731 734 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=136120 $D=0
M2332 120 732 735 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=140750 $D=0
M2333 121 733 736 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=145380 $D=0
M2334 737 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=136120 $D=0
M2335 738 122 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=140750 $D=0
M2336 739 122 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=145380 $D=0
M2337 740 122 115 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=136120 $D=0
M2338 741 122 116 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=140750 $D=0
M2339 742 122 117 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=145380 $D=0
M2340 1045 737 740 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=136120 $D=0
M2341 1046 738 741 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=140750 $D=0
M2342 1047 739 742 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=145380 $D=0
M2343 167 115 1045 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=136120 $D=0
M2344 171 116 1046 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=140750 $D=0
M2345 172 117 1047 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=145380 $D=0
M2346 743 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=136120 $D=0
M2347 744 123 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=140750 $D=0
M2348 745 123 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=145380 $D=0
M2349 124 123 740 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=136120 $D=0
M2350 125 123 741 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=140750 $D=0
M2351 126 123 742 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=145380 $D=0
M2352 11 743 124 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=136120 $D=0
M2353 12 744 125 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=140750 $D=0
M2354 13 745 126 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=145380 $D=0
M2355 748 746 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=136120 $D=0
M2356 749 747 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=140750 $D=0
M2357 750 127 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=145380 $D=0
M2358 167 754 751 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=136120 $D=0
M2359 171 755 752 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=140750 $D=0
M2360 172 756 753 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=145380 $D=0
M2361 757 734 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=136120 $D=0
M2362 758 735 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=140750 $D=0
M2363 759 736 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=145380 $D=0
M2364 754 734 746 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=136120 $D=0
M2365 755 735 747 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=140750 $D=0
M2366 756 736 127 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=145380 $D=0
M2367 748 757 754 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=136120 $D=0
M2368 749 758 755 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=140750 $D=0
M2369 750 759 756 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=145380 $D=0
M2370 760 751 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=136120 $D=0
M2371 761 752 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=140750 $D=0
M2372 762 753 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=145380 $D=0
M2373 128 751 124 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=136120 $D=0
M2374 746 752 125 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=140750 $D=0
M2375 747 753 126 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=145380 $D=0
M2376 734 760 128 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=136120 $D=0
M2377 735 761 746 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=140750 $D=0
M2378 736 762 747 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=145380 $D=0
M2379 763 128 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=136120 $D=0
M2380 764 746 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=140750 $D=0
M2381 765 747 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=145380 $D=0
M2382 766 751 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=136120 $D=0
M2383 767 752 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=140750 $D=0
M2384 768 753 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=145380 $D=0
M2385 769 751 763 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=136120 $D=0
M2386 770 752 764 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=140750 $D=0
M2387 771 753 765 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=145380 $D=0
M2388 124 766 769 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=136120 $D=0
M2389 125 767 770 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=140750 $D=0
M2390 126 768 771 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=145380 $D=0
M2391 1063 734 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=135760 $D=0
M2392 1064 735 171 171 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=140390 $D=0
M2393 1065 736 172 172 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=145020 $D=0
M2394 772 124 1063 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=135760 $D=0
M2395 773 125 1064 171 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=140390 $D=0
M2396 774 126 1065 172 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=145020 $D=0
M2397 775 769 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=136120 $D=0
M2398 776 770 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=140750 $D=0
M2399 777 771 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=145380 $D=0
M2400 778 734 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=136120 $D=0
M2401 779 735 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=140750 $D=0
M2402 780 736 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=145380 $D=0
M2403 167 124 778 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=136120 $D=0
M2404 171 125 779 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=140750 $D=0
M2405 172 126 780 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=145380 $D=0
M2406 781 734 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=136120 $D=0
M2407 782 735 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=140750 $D=0
M2408 783 736 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=145380 $D=0
M2409 167 124 781 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=136120 $D=0
M2410 171 125 782 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=140750 $D=0
M2411 172 126 783 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=145380 $D=0
M2412 1066 734 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=135940 $D=0
M2413 1067 735 171 171 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=140570 $D=0
M2414 1068 736 172 172 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=145200 $D=0
M2415 787 124 1066 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=135940 $D=0
M2416 788 125 1067 171 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=140570 $D=0
M2417 789 126 1068 172 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=145200 $D=0
M2418 167 781 787 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=136120 $D=0
M2419 171 782 788 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=140750 $D=0
M2420 172 783 789 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=145380 $D=0
M2421 790 135 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=136120 $D=0
M2422 791 135 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=140750 $D=0
M2423 792 135 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=145380 $D=0
M2424 793 135 772 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=136120 $D=0
M2425 794 135 773 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=140750 $D=0
M2426 795 135 774 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=145380 $D=0
M2427 778 790 793 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=136120 $D=0
M2428 779 791 794 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=140750 $D=0
M2429 780 792 795 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=145380 $D=0
M2430 796 135 775 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=136120 $D=0
M2431 797 135 776 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=140750 $D=0
M2432 798 135 777 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=145380 $D=0
M2433 787 790 796 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=136120 $D=0
M2434 788 791 797 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=140750 $D=0
M2435 789 792 798 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=145380 $D=0
M2436 799 136 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=136120 $D=0
M2437 800 136 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=140750 $D=0
M2438 801 136 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=145380 $D=0
M2439 802 136 796 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=136120 $D=0
M2440 803 136 797 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=140750 $D=0
M2441 804 136 798 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=145380 $D=0
M2442 793 799 802 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=136120 $D=0
M2443 794 800 803 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=140750 $D=0
M2444 795 801 804 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=145380 $D=0
M2445 14 802 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=136120 $D=0
M2446 15 803 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=140750 $D=0
M2447 16 804 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=145380 $D=0
M2448 805 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=136120 $D=0
M2449 806 137 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=140750 $D=0
M2450 807 137 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=145380 $D=0
M2451 808 137 138 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=136120 $D=0
M2452 809 137 139 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=140750 $D=0
M2453 810 137 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=145380 $D=0
M2454 141 805 808 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=136120 $D=0
M2455 142 806 809 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=140750 $D=0
M2456 138 807 810 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=145380 $D=0
M2457 811 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=136120 $D=0
M2458 812 137 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=140750 $D=0
M2459 813 137 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=145380 $D=0
M2460 814 137 143 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=136120 $D=0
M2461 815 137 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=140750 $D=0
M2462 816 137 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=145380 $D=0
M2463 144 811 814 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=136120 $D=0
M2464 145 812 815 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=140750 $D=0
M2465 146 813 816 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=145380 $D=0
M2466 817 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=136120 $D=0
M2467 818 137 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=140750 $D=0
M2468 819 137 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=145380 $D=0
M2469 820 137 8 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=136120 $D=0
M2470 821 137 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=140750 $D=0
M2471 822 137 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=145380 $D=0
M2472 147 817 820 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=136120 $D=0
M2473 148 818 821 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=140750 $D=0
M2474 149 819 822 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=145380 $D=0
M2475 823 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=136120 $D=0
M2476 824 137 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=140750 $D=0
M2477 825 137 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=145380 $D=0
M2478 826 137 8 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=136120 $D=0
M2479 827 137 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=140750 $D=0
M2480 828 137 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=145380 $D=0
M2481 150 823 826 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=136120 $D=0
M2482 151 824 827 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=140750 $D=0
M2483 152 825 828 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=145380 $D=0
M2484 829 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=136120 $D=0
M2485 830 137 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=140750 $D=0
M2486 831 137 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=145380 $D=0
M2487 832 137 8 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=136120 $D=0
M2488 833 137 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=140750 $D=0
M2489 834 137 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=145380 $D=0
M2490 153 829 832 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=136120 $D=0
M2491 154 830 833 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=140750 $D=0
M2492 155 831 834 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=145380 $D=0
M2493 167 734 1048 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=136120 $D=0
M2494 171 735 1049 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=140750 $D=0
M2495 172 736 1050 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=145380 $D=0
M2496 142 1048 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=136120 $D=0
M2497 138 1049 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=140750 $D=0
M2498 139 1050 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=145380 $D=0
M2499 835 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=136120 $D=0
M2500 836 126 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=140750 $D=0
M2501 837 126 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=145380 $D=0
M2502 146 126 142 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=136120 $D=0
M2503 156 126 138 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=140750 $D=0
M2504 143 126 139 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=145380 $D=0
M2505 808 835 146 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=136120 $D=0
M2506 809 836 156 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=140750 $D=0
M2507 810 837 143 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=145380 $D=0
M2508 838 125 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=136120 $D=0
M2509 839 125 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=140750 $D=0
M2510 840 125 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=145380 $D=0
M2511 134 125 146 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=136120 $D=0
M2512 133 125 156 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=140750 $D=0
M2513 132 125 143 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=145380 $D=0
M2514 814 838 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=136120 $D=0
M2515 815 839 133 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=140750 $D=0
M2516 816 840 132 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=145380 $D=0
M2517 841 124 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=136120 $D=0
M2518 842 124 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=140750 $D=0
M2519 843 124 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=145380 $D=0
M2520 129 124 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=136120 $D=0
M2521 130 124 133 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=140750 $D=0
M2522 131 124 132 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=145380 $D=0
M2523 820 841 129 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=136120 $D=0
M2524 821 842 130 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=140750 $D=0
M2525 822 843 131 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=145380 $D=0
M2526 844 157 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=136120 $D=0
M2527 845 157 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=140750 $D=0
M2528 846 157 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=145380 $D=0
M2529 158 157 129 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=136120 $D=0
M2530 159 157 130 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=140750 $D=0
M2531 160 157 131 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=145380 $D=0
M2532 826 844 158 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=136120 $D=0
M2533 827 845 159 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=140750 $D=0
M2534 828 846 160 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=145380 $D=0
M2535 847 161 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=136120 $D=0
M2536 848 161 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=140750 $D=0
M2537 849 161 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=145380 $D=0
M2538 209 161 158 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=136120 $D=0
M2539 210 161 159 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=140750 $D=0
M2540 211 161 160 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=145380 $D=0
M2541 832 847 209 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=136120 $D=0
M2542 833 848 210 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=140750 $D=0
M2543 834 849 211 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=145380 $D=0
M2544 850 162 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=136120 $D=0
M2545 851 162 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=140750 $D=0
M2546 852 162 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=145380 $D=0
M2547 853 162 115 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=136120 $D=0
M2548 854 162 116 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=140750 $D=0
M2549 855 162 117 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=145380 $D=0
M2550 11 850 853 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=136120 $D=0
M2551 12 851 854 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=140750 $D=0
M2552 13 852 855 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=145380 $D=0
M2553 856 719 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=136120 $D=0
M2554 857 720 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=140750 $D=0
M2555 858 721 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=145380 $D=0
M2556 167 853 856 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=136120 $D=0
M2557 171 854 857 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=140750 $D=0
M2558 172 855 858 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=145380 $D=0
M2559 1069 719 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=135940 $D=0
M2560 1070 720 171 171 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=140570 $D=0
M2561 1071 721 172 172 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=145200 $D=0
M2562 862 853 1069 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=135940 $D=0
M2563 863 854 1070 171 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=140570 $D=0
M2564 864 855 1071 172 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=145200 $D=0
M2565 167 856 862 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=136120 $D=0
M2566 171 857 863 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=140750 $D=0
M2567 172 858 864 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=145380 $D=0
M2568 1051 163 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=136120 $D=0
M2569 1052 865 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=140750 $D=0
M2570 1053 866 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=145380 $D=0
M2571 167 862 1051 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=136120 $D=0
M2572 171 863 1052 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=140750 $D=0
M2573 172 864 1053 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=145380 $D=0
M2574 865 1051 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=136120 $D=0
M2575 866 1052 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=140750 $D=0
M2576 164 1053 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=145380 $D=0
M2577 1072 719 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=135760 $D=0
M2578 1073 720 171 171 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=140390 $D=0
M2579 1074 721 172 172 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=145020 $D=0
M2580 867 870 1072 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=135760 $D=0
M2581 868 871 1073 171 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=140390 $D=0
M2582 869 872 1074 172 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=145020 $D=0
M2583 870 853 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=136120 $D=0
M2584 871 854 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=140750 $D=0
M2585 872 855 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=145380 $D=0
M2586 873 867 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=136120 $D=0
M2587 874 868 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=140750 $D=0
M2588 875 869 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=145380 $D=0
M2589 167 163 873 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=136120 $D=0
M2590 171 865 874 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=140750 $D=0
M2591 172 866 875 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=145380 $D=0
M2592 878 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=136120 $D=0
M2593 879 876 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=140750 $D=0
M2594 880 877 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=145380 $D=0
M2595 876 873 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=136120 $D=0
M2596 877 874 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=140750 $D=0
M2597 166 875 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=145380 $D=0
M2598 167 878 876 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=136120 $D=0
M2599 171 879 877 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=140750 $D=0
M2600 172 880 166 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=145380 $D=0
M2601 883 881 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=136120 $D=0
M2602 884 882 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=140750 $D=0
M2603 885 140 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=145380 $D=0
M2604 167 889 886 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=136120 $D=0
M2605 171 890 887 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=140750 $D=0
M2606 172 891 888 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=145380 $D=0
M2607 892 119 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=136120 $D=0
M2608 893 120 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=140750 $D=0
M2609 894 121 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=145380 $D=0
M2610 889 119 881 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=136120 $D=0
M2611 890 120 882 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=140750 $D=0
M2612 891 121 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=145380 $D=0
M2613 883 892 889 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=136120 $D=0
M2614 884 893 890 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=140750 $D=0
M2615 885 894 891 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=145380 $D=0
M2616 895 886 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=136120 $D=0
M2617 896 887 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=140750 $D=0
M2618 897 888 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=145380 $D=0
M2619 168 886 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=136120 $D=0
M2620 881 887 9 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=140750 $D=0
M2621 882 888 140 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=145380 $D=0
M2622 119 895 168 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=136120 $D=0
M2623 120 896 881 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=140750 $D=0
M2624 121 897 882 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=145380 $D=0
M2625 898 168 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=136120 $D=0
M2626 899 881 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=140750 $D=0
M2627 900 882 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=145380 $D=0
M2628 901 886 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=136120 $D=0
M2629 902 887 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=140750 $D=0
M2630 903 888 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=145380 $D=0
M2631 212 886 898 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=136120 $D=0
M2632 213 887 899 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=140750 $D=0
M2633 214 888 900 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=145380 $D=0
M2634 167 901 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=136120 $D=0
M2635 9 902 213 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=140750 $D=0
M2636 140 903 214 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=145380 $D=0
M2637 904 169 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=136120 $D=0
M2638 905 169 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=140750 $D=0
M2639 906 169 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=145380 $D=0
M2640 907 169 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=136120 $D=0
M2641 908 169 213 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=140750 $D=0
M2642 909 169 214 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=145380 $D=0
M2643 14 904 907 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=136120 $D=0
M2644 15 905 908 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=140750 $D=0
M2645 16 906 909 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=145380 $D=0
M2646 910 170 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=136120 $D=0
M2647 911 170 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=140750 $D=0
M2648 912 170 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=145380 $D=0
M2649 170 170 907 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=136120 $D=0
M2650 170 170 908 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=140750 $D=0
M2651 170 170 909 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=145380 $D=0
M2652 8 910 170 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=136120 $D=0
M2653 9 911 170 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=140750 $D=0
M2654 140 912 170 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=145380 $D=0
M2655 913 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=136120 $D=0
M2656 914 114 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=140750 $D=0
M2657 915 114 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=145380 $D=0
M2658 167 913 916 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=136120 $D=0
M2659 171 914 917 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=140750 $D=0
M2660 172 915 918 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=145380 $D=0
M2661 919 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=136120 $D=0
M2662 920 114 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=140750 $D=0
M2663 921 114 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=145380 $D=0
M2664 922 916 170 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=136120 $D=0
M2665 923 917 170 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=140750 $D=0
M2666 924 918 170 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=145380 $D=0
M2667 167 922 1054 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=136120 $D=0
M2668 171 923 1055 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=140750 $D=0
M2669 172 924 1056 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=145380 $D=0
M2670 925 1054 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=136120 $D=0
M2671 926 1055 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=140750 $D=0
M2672 927 1056 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=145380 $D=0
M2673 922 913 925 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=136120 $D=0
M2674 923 914 926 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=140750 $D=0
M2675 924 915 927 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=145380 $D=0
M2676 928 919 925 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=136120 $D=0
M2677 929 920 926 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=140750 $D=0
M2678 930 921 927 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=145380 $D=0
M2679 167 934 931 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=136120 $D=0
M2680 171 935 932 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=140750 $D=0
M2681 172 936 933 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=145380 $D=0
M2682 934 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=136120 $D=0
M2683 935 114 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=140750 $D=0
M2684 936 114 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=145380 $D=0
M2685 1057 928 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=136120 $D=0
M2686 1058 929 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=140750 $D=0
M2687 1059 930 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=145380 $D=0
M2688 937 934 1057 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=136120 $D=0
M2689 938 935 1058 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=140750 $D=0
M2690 939 936 1059 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=145380 $D=0
M2691 167 937 119 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=136120 $D=0
M2692 171 938 120 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=140750 $D=0
M2693 172 939 121 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=145380 $D=0
M2694 1060 119 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=136120 $D=0
M2695 1061 120 171 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=140750 $D=0
M2696 1062 121 172 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=145380 $D=0
M2697 937 931 1060 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=136120 $D=0
M2698 938 932 1061 171 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=140750 $D=0
M2699 939 933 1062 172 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=145380 $D=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162
** N=788 EP=161 IP=1514 FDC=1800
M0 178 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=125610 $D=1
M1 179 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=130240 $D=1
M2 180 178 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=125610 $D=1
M3 181 179 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=130240 $D=1
M4 7 1 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=125610 $D=1
M5 8 1 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=130240 $D=1
M6 182 178 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=125610 $D=1
M7 183 179 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=130240 $D=1
M8 2 1 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=125610 $D=1
M9 3 1 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=130240 $D=1
M10 184 178 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=125610 $D=1
M11 185 179 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=130240 $D=1
M12 2 1 184 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=125610 $D=1
M13 3 1 185 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=130240 $D=1
M14 188 186 184 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=125610 $D=1
M15 189 187 185 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=130240 $D=1
M16 186 4 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=125610 $D=1
M17 187 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=130240 $D=1
M18 190 186 182 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=125610 $D=1
M19 191 187 183 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=130240 $D=1
M20 180 4 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=125610 $D=1
M21 181 4 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=130240 $D=1
M22 192 5 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=125610 $D=1
M23 193 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=130240 $D=1
M24 194 192 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=125610 $D=1
M25 195 193 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=130240 $D=1
M26 188 5 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=125610 $D=1
M27 189 5 195 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=130240 $D=1
M28 196 6 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=125610 $D=1
M29 197 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=130240 $D=1
M30 198 196 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=125610 $D=1
M31 199 197 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=130240 $D=1
M32 9 6 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=125610 $D=1
M33 10 6 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=130240 $D=1
M34 200 196 11 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=125610 $D=1
M35 201 197 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=130240 $D=1
M36 202 6 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=125610 $D=1
M37 203 6 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=130240 $D=1
M38 206 196 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=125610 $D=1
M39 207 197 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=130240 $D=1
M40 194 6 206 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=125610 $D=1
M41 195 6 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=130240 $D=1
M42 210 208 206 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=125610 $D=1
M43 211 209 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=130240 $D=1
M44 208 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=125610 $D=1
M45 209 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=130240 $D=1
M46 212 208 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=125610 $D=1
M47 213 209 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=130240 $D=1
M48 198 13 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=125610 $D=1
M49 199 13 213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=130240 $D=1
M50 214 14 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=125610 $D=1
M51 215 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=130240 $D=1
M52 216 214 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=125610 $D=1
M53 217 215 213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=130240 $D=1
M54 210 14 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=125610 $D=1
M55 211 14 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=130240 $D=1
M56 7 15 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=125610 $D=1
M57 8 15 219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=130240 $D=1
M58 220 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=125610 $D=1
M59 221 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=130240 $D=1
M60 222 15 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=125610 $D=1
M61 223 15 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=130240 $D=1
M62 7 222 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=125610 $D=1
M63 8 223 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=130240 $D=1
M64 224 687 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=125610 $D=1
M65 225 688 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=130240 $D=1
M66 222 218 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=125610 $D=1
M67 223 219 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=130240 $D=1
M68 224 16 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=125610 $D=1
M69 225 16 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=130240 $D=1
M70 230 17 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=125610 $D=1
M71 231 17 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=130240 $D=1
M72 228 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=125610 $D=1
M73 229 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=130240 $D=1
M74 7 18 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=125610 $D=1
M75 8 18 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=130240 $D=1
M76 234 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=125610 $D=1
M77 235 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=130240 $D=1
M78 236 18 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=125610 $D=1
M79 237 18 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=130240 $D=1
M80 7 236 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=125610 $D=1
M81 8 237 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=130240 $D=1
M82 238 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=125610 $D=1
M83 239 690 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=130240 $D=1
M84 236 232 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=125610 $D=1
M85 237 233 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=130240 $D=1
M86 238 19 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=125610 $D=1
M87 239 19 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=130240 $D=1
M88 230 20 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=125610 $D=1
M89 231 20 239 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=130240 $D=1
M90 240 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=125610 $D=1
M91 241 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=130240 $D=1
M92 7 21 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=125610 $D=1
M93 8 21 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=130240 $D=1
M94 244 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=125610 $D=1
M95 245 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=130240 $D=1
M96 246 21 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=125610 $D=1
M97 247 21 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=130240 $D=1
M98 7 246 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=125610 $D=1
M99 8 247 692 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=130240 $D=1
M100 248 691 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=125610 $D=1
M101 249 692 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=130240 $D=1
M102 246 242 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=125610 $D=1
M103 247 243 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=130240 $D=1
M104 248 22 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=125610 $D=1
M105 249 22 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=130240 $D=1
M106 230 23 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=125610 $D=1
M107 231 23 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=130240 $D=1
M108 250 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=125610 $D=1
M109 251 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=130240 $D=1
M110 7 24 252 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=125610 $D=1
M111 8 24 253 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=130240 $D=1
M112 254 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=125610 $D=1
M113 255 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=130240 $D=1
M114 256 24 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=125610 $D=1
M115 257 24 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=130240 $D=1
M116 7 256 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=125610 $D=1
M117 8 257 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=130240 $D=1
M118 258 693 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=125610 $D=1
M119 259 694 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=130240 $D=1
M120 256 252 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=125610 $D=1
M121 257 253 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=130240 $D=1
M122 258 25 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=125610 $D=1
M123 259 25 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=130240 $D=1
M124 230 26 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=125610 $D=1
M125 231 26 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=130240 $D=1
M126 260 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=125610 $D=1
M127 261 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=130240 $D=1
M128 7 27 262 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=125610 $D=1
M129 8 27 263 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=130240 $D=1
M130 264 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=125610 $D=1
M131 265 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=130240 $D=1
M132 266 27 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=125610 $D=1
M133 267 27 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=130240 $D=1
M134 7 266 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=125610 $D=1
M135 8 267 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=130240 $D=1
M136 268 695 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=125610 $D=1
M137 269 696 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=130240 $D=1
M138 266 262 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=125610 $D=1
M139 267 263 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=130240 $D=1
M140 268 28 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=125610 $D=1
M141 269 28 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=130240 $D=1
M142 230 29 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=125610 $D=1
M143 231 29 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=130240 $D=1
M144 270 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=125610 $D=1
M145 271 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=130240 $D=1
M146 7 30 272 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=125610 $D=1
M147 8 30 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=130240 $D=1
M148 274 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=125610 $D=1
M149 275 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=130240 $D=1
M150 276 30 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=125610 $D=1
M151 277 30 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=130240 $D=1
M152 7 276 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=125610 $D=1
M153 8 277 698 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=130240 $D=1
M154 278 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=125610 $D=1
M155 279 698 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=130240 $D=1
M156 276 272 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=125610 $D=1
M157 277 273 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=130240 $D=1
M158 278 31 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=125610 $D=1
M159 279 31 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=130240 $D=1
M160 230 32 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=125610 $D=1
M161 231 32 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=130240 $D=1
M162 280 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=125610 $D=1
M163 281 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=130240 $D=1
M164 7 33 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=125610 $D=1
M165 8 33 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=130240 $D=1
M166 284 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=125610 $D=1
M167 285 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=130240 $D=1
M168 286 33 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=125610 $D=1
M169 287 33 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=130240 $D=1
M170 7 286 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=125610 $D=1
M171 8 287 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=130240 $D=1
M172 288 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=125610 $D=1
M173 289 700 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=130240 $D=1
M174 286 282 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=125610 $D=1
M175 287 283 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=130240 $D=1
M176 288 34 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=125610 $D=1
M177 289 34 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=130240 $D=1
M178 230 35 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=125610 $D=1
M179 231 35 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=130240 $D=1
M180 290 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=125610 $D=1
M181 291 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=130240 $D=1
M182 7 36 292 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=125610 $D=1
M183 8 36 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=130240 $D=1
M184 294 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=125610 $D=1
M185 295 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=130240 $D=1
M186 296 36 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=125610 $D=1
M187 297 36 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=130240 $D=1
M188 7 296 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=125610 $D=1
M189 8 297 702 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=130240 $D=1
M190 298 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=125610 $D=1
M191 299 702 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=130240 $D=1
M192 296 292 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=125610 $D=1
M193 297 293 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=130240 $D=1
M194 298 37 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=125610 $D=1
M195 299 37 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=130240 $D=1
M196 230 38 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=125610 $D=1
M197 231 38 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=130240 $D=1
M198 300 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=125610 $D=1
M199 301 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=130240 $D=1
M200 7 39 302 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=125610 $D=1
M201 8 39 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=130240 $D=1
M202 304 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=125610 $D=1
M203 305 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=130240 $D=1
M204 306 39 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=125610 $D=1
M205 307 39 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=130240 $D=1
M206 7 306 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=125610 $D=1
M207 8 307 704 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=130240 $D=1
M208 308 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=125610 $D=1
M209 309 704 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=130240 $D=1
M210 306 302 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=125610 $D=1
M211 307 303 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=130240 $D=1
M212 308 40 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=125610 $D=1
M213 309 40 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=130240 $D=1
M214 230 41 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=125610 $D=1
M215 231 41 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=130240 $D=1
M216 310 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=125610 $D=1
M217 311 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=130240 $D=1
M218 7 42 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=125610 $D=1
M219 8 42 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=130240 $D=1
M220 314 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=125610 $D=1
M221 315 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=130240 $D=1
M222 316 42 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=125610 $D=1
M223 317 42 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=130240 $D=1
M224 7 316 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=125610 $D=1
M225 8 317 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=130240 $D=1
M226 318 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=125610 $D=1
M227 319 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=130240 $D=1
M228 316 312 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=125610 $D=1
M229 317 313 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=130240 $D=1
M230 318 43 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=125610 $D=1
M231 319 43 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=130240 $D=1
M232 230 44 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=125610 $D=1
M233 231 44 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=130240 $D=1
M234 320 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=125610 $D=1
M235 321 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=130240 $D=1
M236 7 45 322 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=125610 $D=1
M237 8 45 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=130240 $D=1
M238 324 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=125610 $D=1
M239 325 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=130240 $D=1
M240 326 45 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=125610 $D=1
M241 327 45 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=130240 $D=1
M242 7 326 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=125610 $D=1
M243 8 327 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=130240 $D=1
M244 328 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=125610 $D=1
M245 329 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=130240 $D=1
M246 326 322 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=125610 $D=1
M247 327 323 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=130240 $D=1
M248 328 46 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=125610 $D=1
M249 329 46 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=130240 $D=1
M250 230 47 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=125610 $D=1
M251 231 47 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=130240 $D=1
M252 330 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=125610 $D=1
M253 331 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=130240 $D=1
M254 7 48 332 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=125610 $D=1
M255 8 48 333 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=130240 $D=1
M256 334 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=125610 $D=1
M257 335 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=130240 $D=1
M258 336 48 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=125610 $D=1
M259 337 48 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=130240 $D=1
M260 7 336 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=125610 $D=1
M261 8 337 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=130240 $D=1
M262 338 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=125610 $D=1
M263 339 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=130240 $D=1
M264 336 332 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=125610 $D=1
M265 337 333 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=130240 $D=1
M266 338 49 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=125610 $D=1
M267 339 49 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=130240 $D=1
M268 230 50 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=125610 $D=1
M269 231 50 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=130240 $D=1
M270 340 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=125610 $D=1
M271 341 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=130240 $D=1
M272 7 51 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=125610 $D=1
M273 8 51 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=130240 $D=1
M274 344 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=125610 $D=1
M275 345 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=130240 $D=1
M276 346 51 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=125610 $D=1
M277 347 51 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=130240 $D=1
M278 7 346 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=125610 $D=1
M279 8 347 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=130240 $D=1
M280 348 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=125610 $D=1
M281 349 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=130240 $D=1
M282 346 342 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=125610 $D=1
M283 347 343 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=130240 $D=1
M284 348 52 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=125610 $D=1
M285 349 52 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=130240 $D=1
M286 230 53 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=125610 $D=1
M287 231 53 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=130240 $D=1
M288 350 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=125610 $D=1
M289 351 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=130240 $D=1
M290 7 54 352 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=125610 $D=1
M291 8 54 353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=130240 $D=1
M292 354 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=125610 $D=1
M293 355 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=130240 $D=1
M294 356 54 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=125610 $D=1
M295 357 54 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=130240 $D=1
M296 7 356 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=125610 $D=1
M297 8 357 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=130240 $D=1
M298 358 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=125610 $D=1
M299 359 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=130240 $D=1
M300 356 352 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=125610 $D=1
M301 357 353 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=130240 $D=1
M302 358 55 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=125610 $D=1
M303 359 55 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=130240 $D=1
M304 230 56 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=125610 $D=1
M305 231 56 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=130240 $D=1
M306 360 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=125610 $D=1
M307 361 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=130240 $D=1
M308 7 57 362 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=125610 $D=1
M309 8 57 363 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=130240 $D=1
M310 364 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=125610 $D=1
M311 365 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=130240 $D=1
M312 366 57 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=125610 $D=1
M313 367 57 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=130240 $D=1
M314 7 366 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=125610 $D=1
M315 8 367 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=130240 $D=1
M316 368 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=125610 $D=1
M317 369 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=130240 $D=1
M318 366 362 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=125610 $D=1
M319 367 363 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=130240 $D=1
M320 368 58 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=125610 $D=1
M321 369 58 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=130240 $D=1
M322 230 59 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=125610 $D=1
M323 231 59 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=130240 $D=1
M324 370 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=125610 $D=1
M325 371 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=130240 $D=1
M326 7 60 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=125610 $D=1
M327 8 60 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=130240 $D=1
M328 374 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=125610 $D=1
M329 375 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=130240 $D=1
M330 376 60 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=125610 $D=1
M331 377 60 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=130240 $D=1
M332 7 376 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=125610 $D=1
M333 8 377 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=130240 $D=1
M334 378 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=125610 $D=1
M335 379 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=130240 $D=1
M336 376 372 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=125610 $D=1
M337 377 373 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=130240 $D=1
M338 378 61 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=125610 $D=1
M339 379 61 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=130240 $D=1
M340 230 62 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=125610 $D=1
M341 231 62 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=130240 $D=1
M342 380 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=125610 $D=1
M343 381 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=130240 $D=1
M344 7 63 382 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=125610 $D=1
M345 8 63 383 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=130240 $D=1
M346 384 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=125610 $D=1
M347 385 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=130240 $D=1
M348 386 63 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=125610 $D=1
M349 387 63 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=130240 $D=1
M350 7 386 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=125610 $D=1
M351 8 387 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=130240 $D=1
M352 388 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=125610 $D=1
M353 389 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=130240 $D=1
M354 386 382 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=125610 $D=1
M355 387 383 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=130240 $D=1
M356 388 64 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=125610 $D=1
M357 389 64 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=130240 $D=1
M358 230 65 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=125610 $D=1
M359 231 65 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=130240 $D=1
M360 390 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=125610 $D=1
M361 391 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=130240 $D=1
M362 7 66 392 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=125610 $D=1
M363 8 66 393 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=130240 $D=1
M364 394 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=125610 $D=1
M365 395 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=130240 $D=1
M366 396 66 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=125610 $D=1
M367 397 66 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=130240 $D=1
M368 7 396 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=125610 $D=1
M369 8 397 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=130240 $D=1
M370 398 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=125610 $D=1
M371 399 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=130240 $D=1
M372 396 392 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=125610 $D=1
M373 397 393 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=130240 $D=1
M374 398 67 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=125610 $D=1
M375 399 67 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=130240 $D=1
M376 230 68 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=125610 $D=1
M377 231 68 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=130240 $D=1
M378 400 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=125610 $D=1
M379 401 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=130240 $D=1
M380 7 69 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=125610 $D=1
M381 8 69 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=130240 $D=1
M382 404 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=125610 $D=1
M383 405 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=130240 $D=1
M384 406 69 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=125610 $D=1
M385 407 69 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=130240 $D=1
M386 7 406 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=125610 $D=1
M387 8 407 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=130240 $D=1
M388 408 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=125610 $D=1
M389 409 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=130240 $D=1
M390 406 402 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=125610 $D=1
M391 407 403 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=130240 $D=1
M392 408 70 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=125610 $D=1
M393 409 70 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=130240 $D=1
M394 230 71 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=125610 $D=1
M395 231 71 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=130240 $D=1
M396 410 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=125610 $D=1
M397 411 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=130240 $D=1
M398 7 72 412 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=125610 $D=1
M399 8 72 413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=130240 $D=1
M400 414 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=125610 $D=1
M401 415 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=130240 $D=1
M402 416 72 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=125610 $D=1
M403 417 72 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=130240 $D=1
M404 7 416 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=125610 $D=1
M405 8 417 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=130240 $D=1
M406 418 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=125610 $D=1
M407 419 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=130240 $D=1
M408 416 412 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=125610 $D=1
M409 417 413 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=130240 $D=1
M410 418 73 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=125610 $D=1
M411 419 73 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=130240 $D=1
M412 230 74 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=125610 $D=1
M413 231 74 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=130240 $D=1
M414 420 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=125610 $D=1
M415 421 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=130240 $D=1
M416 7 75 422 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=125610 $D=1
M417 8 75 423 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=130240 $D=1
M418 424 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=125610 $D=1
M419 425 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=130240 $D=1
M420 426 75 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=125610 $D=1
M421 427 75 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=130240 $D=1
M422 7 426 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=125610 $D=1
M423 8 427 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=130240 $D=1
M424 428 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=125610 $D=1
M425 429 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=130240 $D=1
M426 426 422 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=125610 $D=1
M427 427 423 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=130240 $D=1
M428 428 76 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=125610 $D=1
M429 429 76 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=130240 $D=1
M430 230 77 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=125610 $D=1
M431 231 77 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=130240 $D=1
M432 430 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=125610 $D=1
M433 431 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=130240 $D=1
M434 7 78 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=125610 $D=1
M435 8 78 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=130240 $D=1
M436 434 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=125610 $D=1
M437 435 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=130240 $D=1
M438 436 78 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=125610 $D=1
M439 437 78 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=130240 $D=1
M440 7 436 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=125610 $D=1
M441 8 437 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=130240 $D=1
M442 438 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=125610 $D=1
M443 439 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=130240 $D=1
M444 436 432 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=125610 $D=1
M445 437 433 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=130240 $D=1
M446 438 79 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=125610 $D=1
M447 439 79 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=130240 $D=1
M448 230 80 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=125610 $D=1
M449 231 80 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=130240 $D=1
M450 440 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=125610 $D=1
M451 441 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=130240 $D=1
M452 7 81 442 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=125610 $D=1
M453 8 81 443 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=130240 $D=1
M454 444 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=125610 $D=1
M455 445 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=130240 $D=1
M456 446 81 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=125610 $D=1
M457 447 81 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=130240 $D=1
M458 7 446 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=125610 $D=1
M459 8 447 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=130240 $D=1
M460 448 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=125610 $D=1
M461 449 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=130240 $D=1
M462 446 442 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=125610 $D=1
M463 447 443 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=130240 $D=1
M464 448 82 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=125610 $D=1
M465 449 82 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=130240 $D=1
M466 230 83 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=125610 $D=1
M467 231 83 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=130240 $D=1
M468 450 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=125610 $D=1
M469 451 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=130240 $D=1
M470 7 84 452 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=125610 $D=1
M471 8 84 453 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=130240 $D=1
M472 454 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=125610 $D=1
M473 455 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=130240 $D=1
M474 456 84 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=125610 $D=1
M475 457 84 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=130240 $D=1
M476 7 456 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=125610 $D=1
M477 8 457 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=130240 $D=1
M478 458 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=125610 $D=1
M479 459 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=130240 $D=1
M480 456 452 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=125610 $D=1
M481 457 453 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=130240 $D=1
M482 458 85 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=125610 $D=1
M483 459 85 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=130240 $D=1
M484 230 86 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=125610 $D=1
M485 231 86 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=130240 $D=1
M486 460 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=125610 $D=1
M487 461 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=130240 $D=1
M488 7 87 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=125610 $D=1
M489 8 87 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=130240 $D=1
M490 464 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=125610 $D=1
M491 465 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=130240 $D=1
M492 466 87 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=125610 $D=1
M493 467 87 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=130240 $D=1
M494 7 466 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=125610 $D=1
M495 8 467 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=130240 $D=1
M496 468 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=125610 $D=1
M497 469 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=130240 $D=1
M498 466 462 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=125610 $D=1
M499 467 463 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=130240 $D=1
M500 468 88 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=125610 $D=1
M501 469 88 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=130240 $D=1
M502 230 89 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=125610 $D=1
M503 231 89 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=130240 $D=1
M504 470 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=125610 $D=1
M505 471 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=130240 $D=1
M506 7 90 472 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=125610 $D=1
M507 8 90 473 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=130240 $D=1
M508 474 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=125610 $D=1
M509 475 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=130240 $D=1
M510 476 90 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=125610 $D=1
M511 477 90 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=130240 $D=1
M512 7 476 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=125610 $D=1
M513 8 477 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=130240 $D=1
M514 478 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=125610 $D=1
M515 479 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=130240 $D=1
M516 476 472 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=125610 $D=1
M517 477 473 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=130240 $D=1
M518 478 91 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=125610 $D=1
M519 479 91 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=130240 $D=1
M520 230 92 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=125610 $D=1
M521 231 92 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=130240 $D=1
M522 480 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=125610 $D=1
M523 481 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=130240 $D=1
M524 7 93 482 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=125610 $D=1
M525 8 93 483 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=130240 $D=1
M526 484 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=125610 $D=1
M527 485 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=130240 $D=1
M528 486 93 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=125610 $D=1
M529 487 93 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=130240 $D=1
M530 7 486 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=125610 $D=1
M531 8 487 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=130240 $D=1
M532 488 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=125610 $D=1
M533 489 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=130240 $D=1
M534 486 482 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=125610 $D=1
M535 487 483 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=130240 $D=1
M536 488 94 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=125610 $D=1
M537 489 94 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=130240 $D=1
M538 230 95 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=125610 $D=1
M539 231 95 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=130240 $D=1
M540 490 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=125610 $D=1
M541 491 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=130240 $D=1
M542 7 96 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=125610 $D=1
M543 8 96 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=130240 $D=1
M544 494 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=125610 $D=1
M545 495 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=130240 $D=1
M546 496 96 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=125610 $D=1
M547 497 96 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=130240 $D=1
M548 7 496 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=125610 $D=1
M549 8 497 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=130240 $D=1
M550 498 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=125610 $D=1
M551 499 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=130240 $D=1
M552 496 492 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=125610 $D=1
M553 497 493 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=130240 $D=1
M554 498 97 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=125610 $D=1
M555 499 97 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=130240 $D=1
M556 230 98 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=125610 $D=1
M557 231 98 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=130240 $D=1
M558 500 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=125610 $D=1
M559 501 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=130240 $D=1
M560 7 99 502 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=125610 $D=1
M561 8 99 503 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=130240 $D=1
M562 504 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=125610 $D=1
M563 505 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=130240 $D=1
M564 506 99 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=125610 $D=1
M565 507 99 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=130240 $D=1
M566 7 506 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=125610 $D=1
M567 8 507 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=130240 $D=1
M568 508 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=125610 $D=1
M569 509 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=130240 $D=1
M570 506 502 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=125610 $D=1
M571 507 503 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=130240 $D=1
M572 508 100 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=125610 $D=1
M573 509 100 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=130240 $D=1
M574 230 101 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=125610 $D=1
M575 231 101 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=130240 $D=1
M576 510 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=125610 $D=1
M577 511 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=130240 $D=1
M578 7 102 512 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=125610 $D=1
M579 8 102 513 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=130240 $D=1
M580 514 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=125610 $D=1
M581 515 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=130240 $D=1
M582 516 102 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=125610 $D=1
M583 517 102 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=130240 $D=1
M584 7 516 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=125610 $D=1
M585 8 517 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=130240 $D=1
M586 518 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=125610 $D=1
M587 519 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=130240 $D=1
M588 516 512 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=125610 $D=1
M589 517 513 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=130240 $D=1
M590 518 103 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=125610 $D=1
M591 519 103 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=130240 $D=1
M592 230 104 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=125610 $D=1
M593 231 104 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=130240 $D=1
M594 520 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=125610 $D=1
M595 521 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=130240 $D=1
M596 7 105 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=125610 $D=1
M597 8 105 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=130240 $D=1
M598 524 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=125610 $D=1
M599 525 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=130240 $D=1
M600 526 105 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=125610 $D=1
M601 527 105 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=130240 $D=1
M602 7 526 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=125610 $D=1
M603 8 527 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=130240 $D=1
M604 528 747 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=125610 $D=1
M605 529 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=130240 $D=1
M606 526 522 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=125610 $D=1
M607 527 523 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=130240 $D=1
M608 528 106 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=125610 $D=1
M609 529 106 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=130240 $D=1
M610 230 107 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=125610 $D=1
M611 231 107 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=130240 $D=1
M612 530 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=125610 $D=1
M613 531 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=130240 $D=1
M614 7 108 532 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=125610 $D=1
M615 8 108 533 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=130240 $D=1
M616 534 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=125610 $D=1
M617 535 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=130240 $D=1
M618 7 109 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=125610 $D=1
M619 8 109 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=130240 $D=1
M620 230 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=125610 $D=1
M621 231 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=130240 $D=1
M622 7 538 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=125610 $D=1
M623 8 539 537 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=130240 $D=1
M624 538 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=125610 $D=1
M625 539 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=130240 $D=1
M626 749 226 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=125610 $D=1
M627 750 227 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=130240 $D=1
M628 540 536 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=125610 $D=1
M629 541 537 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=130240 $D=1
M630 7 540 542 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=125610 $D=1
M631 8 541 543 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=130240 $D=1
M632 751 542 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=125610 $D=1
M633 752 543 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=130240 $D=1
M634 540 538 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=125610 $D=1
M635 541 539 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=130240 $D=1
M636 7 546 544 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=125610 $D=1
M637 8 547 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=130240 $D=1
M638 546 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=125610 $D=1
M639 547 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=130240 $D=1
M640 753 230 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=125610 $D=1
M641 754 231 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=130240 $D=1
M642 548 544 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=125610 $D=1
M643 549 545 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=130240 $D=1
M644 7 548 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=125610 $D=1
M645 8 549 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=130240 $D=1
M646 755 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=125610 $D=1
M647 756 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=130240 $D=1
M648 548 546 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=125610 $D=1
M649 549 547 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=130240 $D=1
M650 550 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=125610 $D=1
M651 551 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=130240 $D=1
M652 552 550 542 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=125610 $D=1
M653 553 551 543 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=130240 $D=1
M654 114 113 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=125610 $D=1
M655 115 113 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=130240 $D=1
M656 554 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=125610 $D=1
M657 555 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=130240 $D=1
M658 556 554 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=125610 $D=1
M659 557 555 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=130240 $D=1
M660 757 116 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=125610 $D=1
M661 758 116 557 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=130240 $D=1
M662 7 111 757 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=125610 $D=1
M663 8 112 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=130240 $D=1
M664 558 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=125610 $D=1
M665 559 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=130240 $D=1
M666 118 558 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=125610 $D=1
M667 119 559 557 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=130240 $D=1
M668 9 117 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=125610 $D=1
M669 10 117 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=130240 $D=1
M670 561 560 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=125610 $D=1
M671 562 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=130240 $D=1
M672 7 565 563 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=125610 $D=1
M673 8 566 564 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=130240 $D=1
M674 567 552 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=125610 $D=1
M675 568 553 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=130240 $D=1
M676 565 567 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=125610 $D=1
M677 566 568 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=130240 $D=1
M678 561 552 565 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=125610 $D=1
M679 562 553 566 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=130240 $D=1
M680 569 563 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=125610 $D=1
M681 570 564 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=130240 $D=1
M682 571 569 118 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=125610 $D=1
M683 560 570 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=130240 $D=1
M684 552 563 571 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=125610 $D=1
M685 553 564 560 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=130240 $D=1
M686 572 571 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=125610 $D=1
M687 573 560 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=130240 $D=1
M688 574 563 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=125610 $D=1
M689 575 564 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=130240 $D=1
M690 576 574 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=125610 $D=1
M691 577 575 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=130240 $D=1
M692 118 563 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=125610 $D=1
M693 119 564 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=130240 $D=1
M694 578 552 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=125610 $D=1
M695 579 553 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=130240 $D=1
M696 7 118 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=125610 $D=1
M697 8 119 579 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=130240 $D=1
M698 580 576 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=125610 $D=1
M699 581 577 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=130240 $D=1
M700 777 552 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=125610 $D=1
M701 778 553 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=130240 $D=1
M702 582 118 777 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=125610 $D=1
M703 583 119 778 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=130240 $D=1
M704 779 552 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=125610 $D=1
M705 780 553 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=130240 $D=1
M706 584 118 779 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=125610 $D=1
M707 585 119 780 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=130240 $D=1
M708 588 552 586 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=125610 $D=1
M709 589 553 587 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=130240 $D=1
M710 586 118 588 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=125610 $D=1
M711 587 119 589 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=130240 $D=1
M712 7 584 586 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=125610 $D=1
M713 8 585 587 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=130240 $D=1
M714 590 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=125610 $D=1
M715 591 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=130240 $D=1
M716 592 590 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=125610 $D=1
M717 593 591 579 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=130240 $D=1
M718 582 126 592 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=125610 $D=1
M719 583 126 593 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=130240 $D=1
M720 594 590 580 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=125610 $D=1
M721 595 591 581 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=130240 $D=1
M722 588 126 594 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=125610 $D=1
M723 589 126 595 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=130240 $D=1
M724 596 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=125610 $D=1
M725 597 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=130240 $D=1
M726 598 596 594 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=125610 $D=1
M727 599 597 595 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=130240 $D=1
M728 592 127 598 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=125610 $D=1
M729 593 127 599 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=130240 $D=1
M730 11 598 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=125610 $D=1
M731 12 599 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=130240 $D=1
M732 600 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=125610 $D=1
M733 601 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=130240 $D=1
M734 602 600 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=125610 $D=1
M735 603 601 131 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=130240 $D=1
M736 132 129 602 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=125610 $D=1
M737 133 129 603 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=130240 $D=1
M738 604 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=125610 $D=1
M739 605 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=130240 $D=1
M740 606 604 134 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=125610 $D=1
M741 607 605 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=130240 $D=1
M742 136 129 606 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=125610 $D=1
M743 137 129 607 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=130240 $D=1
M744 608 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=125610 $D=1
M745 609 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=130240 $D=1
M746 138 608 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=125610 $D=1
M747 138 609 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=130240 $D=1
M748 128 129 138 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=125610 $D=1
M749 139 129 138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=130240 $D=1
M750 610 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=125610 $D=1
M751 611 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=130240 $D=1
M752 612 610 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=125610 $D=1
M753 613 611 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=130240 $D=1
M754 140 129 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=125610 $D=1
M755 141 129 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=130240 $D=1
M756 614 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=125610 $D=1
M757 615 129 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=130240 $D=1
M758 616 614 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=125610 $D=1
M759 617 615 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=130240 $D=1
M760 142 129 616 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=125610 $D=1
M761 143 129 617 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=130240 $D=1
M762 7 552 759 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=125610 $D=1
M763 8 553 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=130240 $D=1
M764 133 759 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=125610 $D=1
M765 130 760 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=130240 $D=1
M766 618 144 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=125610 $D=1
M767 619 144 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=130240 $D=1
M768 145 618 133 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=125610 $D=1
M769 146 619 130 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=130240 $D=1
M770 602 144 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=125610 $D=1
M771 603 144 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=130240 $D=1
M772 620 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=125610 $D=1
M773 621 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=130240 $D=1
M774 148 620 145 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=125610 $D=1
M775 125 621 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=130240 $D=1
M776 606 147 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=125610 $D=1
M777 607 147 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=130240 $D=1
M778 622 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=125610 $D=1
M779 623 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=130240 $D=1
M780 121 622 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=125610 $D=1
M781 122 623 125 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=130240 $D=1
M782 138 149 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=125610 $D=1
M783 138 149 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=130240 $D=1
M784 624 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=125610 $D=1
M785 625 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=130240 $D=1
M786 150 624 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=125610 $D=1
M787 151 625 122 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=130240 $D=1
M788 612 119 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=125610 $D=1
M789 613 119 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=130240 $D=1
M790 626 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=125610 $D=1
M791 627 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=130240 $D=1
M792 202 626 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=125610 $D=1
M793 203 627 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=130240 $D=1
M794 616 118 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=125610 $D=1
M795 617 118 203 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=130240 $D=1
M796 628 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=125610 $D=1
M797 629 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=130240 $D=1
M798 630 628 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=125610 $D=1
M799 631 629 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=130240 $D=1
M800 9 152 630 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=125610 $D=1
M801 10 152 631 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=130240 $D=1
M802 781 542 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=125610 $D=1
M803 782 543 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=130240 $D=1
M804 632 630 781 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=125610 $D=1
M805 633 631 782 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=130240 $D=1
M806 636 542 634 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=125610 $D=1
M807 637 543 635 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=130240 $D=1
M808 634 630 636 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=125610 $D=1
M809 635 631 637 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=130240 $D=1
M810 7 632 634 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=125610 $D=1
M811 8 633 635 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=130240 $D=1
M812 783 153 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=125610 $D=1
M813 784 638 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=130240 $D=1
M814 761 636 783 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=125610 $D=1
M815 762 637 784 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=130240 $D=1
M816 638 761 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=125610 $D=1
M817 154 762 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=130240 $D=1
M818 639 542 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=125610 $D=1
M819 640 543 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=130240 $D=1
M820 7 641 639 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=125610 $D=1
M821 8 642 640 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=130240 $D=1
M822 641 630 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=125610 $D=1
M823 642 631 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=130240 $D=1
M824 785 639 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=125610 $D=1
M825 786 640 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=130240 $D=1
M826 643 153 785 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=125610 $D=1
M827 644 638 786 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=130240 $D=1
M828 646 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=125610 $D=1
M829 647 645 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=130240 $D=1
M830 787 643 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=125610 $D=1
M831 788 644 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=130240 $D=1
M832 645 646 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=125610 $D=1
M833 156 647 788 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=130240 $D=1
M834 649 648 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=125610 $D=1
M835 650 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=130240 $D=1
M836 7 653 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=125610 $D=1
M837 8 654 652 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=130240 $D=1
M838 655 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=125610 $D=1
M839 656 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=130240 $D=1
M840 653 655 648 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=125610 $D=1
M841 654 656 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=130240 $D=1
M842 649 114 653 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=125610 $D=1
M843 650 115 654 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=130240 $D=1
M844 657 651 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=125610 $D=1
M845 658 652 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=130240 $D=1
M846 158 657 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=125610 $D=1
M847 648 658 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=130240 $D=1
M848 114 651 158 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=125610 $D=1
M849 115 652 648 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=130240 $D=1
M850 659 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=125610 $D=1
M851 660 648 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=130240 $D=1
M852 661 651 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=125610 $D=1
M853 662 652 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=130240 $D=1
M854 204 661 659 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=125610 $D=1
M855 205 662 660 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=130240 $D=1
M856 7 651 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=125610 $D=1
M857 8 652 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=130240 $D=1
M858 663 159 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=125610 $D=1
M859 664 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=130240 $D=1
M860 665 663 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=125610 $D=1
M861 666 664 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=130240 $D=1
M862 11 159 665 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=125610 $D=1
M863 12 159 666 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=130240 $D=1
M864 667 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=125610 $D=1
M865 668 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=130240 $D=1
M866 160 667 665 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=125610 $D=1
M867 160 668 666 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=130240 $D=1
M868 7 160 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=125610 $D=1
M869 8 160 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=130240 $D=1
M870 669 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=125610 $D=1
M871 670 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=130240 $D=1
M872 7 669 671 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=125610 $D=1
M873 8 670 672 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=130240 $D=1
M874 673 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=125610 $D=1
M875 674 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=130240 $D=1
M876 675 669 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=125610 $D=1
M877 676 670 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=130240 $D=1
M878 7 675 763 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=125610 $D=1
M879 8 676 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=130240 $D=1
M880 677 763 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=125610 $D=1
M881 678 764 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=130240 $D=1
M882 675 671 677 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=125610 $D=1
M883 676 672 678 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=130240 $D=1
M884 679 110 677 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=125610 $D=1
M885 680 110 678 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=130240 $D=1
M886 7 683 681 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=125610 $D=1
M887 8 684 682 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=130240 $D=1
M888 683 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=125610 $D=1
M889 684 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=130240 $D=1
M890 765 679 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=125610 $D=1
M891 766 680 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=130240 $D=1
M892 685 681 765 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=125610 $D=1
M893 686 682 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=130240 $D=1
M894 7 685 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=125610 $D=1
M895 8 686 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=130240 $D=1
M896 767 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=125610 $D=1
M897 768 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=130240 $D=1
M898 685 683 767 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=125610 $D=1
M899 686 684 768 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=130240 $D=1
M900 178 1 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=126860 $D=0
M901 179 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=131490 $D=0
M902 180 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=126860 $D=0
M903 181 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=131490 $D=0
M904 7 178 180 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=126860 $D=0
M905 8 179 181 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=131490 $D=0
M906 182 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=126860 $D=0
M907 183 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=131490 $D=0
M908 2 178 182 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=126860 $D=0
M909 3 179 183 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=131490 $D=0
M910 184 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=126860 $D=0
M911 185 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=131490 $D=0
M912 2 178 184 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=126860 $D=0
M913 3 179 185 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=131490 $D=0
M914 188 4 184 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=126860 $D=0
M915 189 4 185 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=131490 $D=0
M916 186 4 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=126860 $D=0
M917 187 4 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=131490 $D=0
M918 190 4 182 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=126860 $D=0
M919 191 4 183 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=131490 $D=0
M920 180 186 190 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=126860 $D=0
M921 181 187 191 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=131490 $D=0
M922 192 5 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=126860 $D=0
M923 193 5 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=131490 $D=0
M924 194 5 190 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=126860 $D=0
M925 195 5 191 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=131490 $D=0
M926 188 192 194 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=126860 $D=0
M927 189 193 195 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=131490 $D=0
M928 196 6 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=126860 $D=0
M929 197 6 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=131490 $D=0
M930 198 6 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=126860 $D=0
M931 199 6 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=131490 $D=0
M932 9 196 198 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=126860 $D=0
M933 10 197 199 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=131490 $D=0
M934 200 6 11 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=126860 $D=0
M935 201 6 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=131490 $D=0
M936 202 196 200 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=126860 $D=0
M937 203 197 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=131490 $D=0
M938 206 6 204 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=126860 $D=0
M939 207 6 205 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=131490 $D=0
M940 194 196 206 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=126860 $D=0
M941 195 197 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=131490 $D=0
M942 210 13 206 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=126860 $D=0
M943 211 13 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=131490 $D=0
M944 208 13 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=126860 $D=0
M945 209 13 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=131490 $D=0
M946 212 13 200 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=126860 $D=0
M947 213 13 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=131490 $D=0
M948 198 208 212 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=126860 $D=0
M949 199 209 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=131490 $D=0
M950 214 14 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=126860 $D=0
M951 215 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=131490 $D=0
M952 216 14 212 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=126860 $D=0
M953 217 14 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=131490 $D=0
M954 210 214 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=126860 $D=0
M955 211 215 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=131490 $D=0
M956 161 15 218 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=126860 $D=0
M957 162 15 219 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=131490 $D=0
M958 220 16 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=126860 $D=0
M959 221 16 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=131490 $D=0
M960 222 218 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=126860 $D=0
M961 223 219 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=131490 $D=0
M962 161 222 687 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=126860 $D=0
M963 162 223 688 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=131490 $D=0
M964 224 687 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=126860 $D=0
M965 225 688 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=131490 $D=0
M966 222 15 224 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=126860 $D=0
M967 223 15 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=131490 $D=0
M968 224 220 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=126860 $D=0
M969 225 221 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=131490 $D=0
M970 230 228 224 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=126860 $D=0
M971 231 229 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=131490 $D=0
M972 228 17 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=126860 $D=0
M973 229 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=131490 $D=0
M974 161 18 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=126860 $D=0
M975 162 18 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=131490 $D=0
M976 234 19 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=126860 $D=0
M977 235 19 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=131490 $D=0
M978 236 232 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=126860 $D=0
M979 237 233 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=131490 $D=0
M980 161 236 689 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=126860 $D=0
M981 162 237 690 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=131490 $D=0
M982 238 689 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=126860 $D=0
M983 239 690 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=131490 $D=0
M984 236 18 238 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=126860 $D=0
M985 237 18 239 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=131490 $D=0
M986 238 234 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=126860 $D=0
M987 239 235 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=131490 $D=0
M988 230 240 238 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=126860 $D=0
M989 231 241 239 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=131490 $D=0
M990 240 20 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=126860 $D=0
M991 241 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=131490 $D=0
M992 161 21 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=126860 $D=0
M993 162 21 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=131490 $D=0
M994 244 22 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=126860 $D=0
M995 245 22 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=131490 $D=0
M996 246 242 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=126860 $D=0
M997 247 243 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=131490 $D=0
M998 161 246 691 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=126860 $D=0
M999 162 247 692 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=131490 $D=0
M1000 248 691 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=126860 $D=0
M1001 249 692 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=131490 $D=0
M1002 246 21 248 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=126860 $D=0
M1003 247 21 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=131490 $D=0
M1004 248 244 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=126860 $D=0
M1005 249 245 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=131490 $D=0
M1006 230 250 248 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=126860 $D=0
M1007 231 251 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=131490 $D=0
M1008 250 23 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=126860 $D=0
M1009 251 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=131490 $D=0
M1010 161 24 252 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=126860 $D=0
M1011 162 24 253 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=131490 $D=0
M1012 254 25 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=126860 $D=0
M1013 255 25 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=131490 $D=0
M1014 256 252 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=126860 $D=0
M1015 257 253 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=131490 $D=0
M1016 161 256 693 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=126860 $D=0
M1017 162 257 694 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=131490 $D=0
M1018 258 693 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=126860 $D=0
M1019 259 694 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=131490 $D=0
M1020 256 24 258 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=126860 $D=0
M1021 257 24 259 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=131490 $D=0
M1022 258 254 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=126860 $D=0
M1023 259 255 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=131490 $D=0
M1024 230 260 258 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=126860 $D=0
M1025 231 261 259 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=131490 $D=0
M1026 260 26 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=126860 $D=0
M1027 261 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=131490 $D=0
M1028 161 27 262 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=126860 $D=0
M1029 162 27 263 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=131490 $D=0
M1030 264 28 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=126860 $D=0
M1031 265 28 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=131490 $D=0
M1032 266 262 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=126860 $D=0
M1033 267 263 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=131490 $D=0
M1034 161 266 695 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=126860 $D=0
M1035 162 267 696 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=131490 $D=0
M1036 268 695 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=126860 $D=0
M1037 269 696 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=131490 $D=0
M1038 266 27 268 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=126860 $D=0
M1039 267 27 269 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=131490 $D=0
M1040 268 264 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=126860 $D=0
M1041 269 265 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=131490 $D=0
M1042 230 270 268 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=126860 $D=0
M1043 231 271 269 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=131490 $D=0
M1044 270 29 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=126860 $D=0
M1045 271 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=131490 $D=0
M1046 161 30 272 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=126860 $D=0
M1047 162 30 273 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=131490 $D=0
M1048 274 31 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=126860 $D=0
M1049 275 31 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=131490 $D=0
M1050 276 272 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=126860 $D=0
M1051 277 273 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=131490 $D=0
M1052 161 276 697 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=126860 $D=0
M1053 162 277 698 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=131490 $D=0
M1054 278 697 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=126860 $D=0
M1055 279 698 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=131490 $D=0
M1056 276 30 278 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=126860 $D=0
M1057 277 30 279 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=131490 $D=0
M1058 278 274 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=126860 $D=0
M1059 279 275 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=131490 $D=0
M1060 230 280 278 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=126860 $D=0
M1061 231 281 279 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=131490 $D=0
M1062 280 32 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=126860 $D=0
M1063 281 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=131490 $D=0
M1064 161 33 282 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=126860 $D=0
M1065 162 33 283 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=131490 $D=0
M1066 284 34 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=126860 $D=0
M1067 285 34 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=131490 $D=0
M1068 286 282 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=126860 $D=0
M1069 287 283 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=131490 $D=0
M1070 161 286 699 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=126860 $D=0
M1071 162 287 700 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=131490 $D=0
M1072 288 699 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=126860 $D=0
M1073 289 700 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=131490 $D=0
M1074 286 33 288 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=126860 $D=0
M1075 287 33 289 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=131490 $D=0
M1076 288 284 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=126860 $D=0
M1077 289 285 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=131490 $D=0
M1078 230 290 288 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=126860 $D=0
M1079 231 291 289 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=131490 $D=0
M1080 290 35 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=126860 $D=0
M1081 291 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=131490 $D=0
M1082 161 36 292 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=126860 $D=0
M1083 162 36 293 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=131490 $D=0
M1084 294 37 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=126860 $D=0
M1085 295 37 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=131490 $D=0
M1086 296 292 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=126860 $D=0
M1087 297 293 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=131490 $D=0
M1088 161 296 701 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=126860 $D=0
M1089 162 297 702 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=131490 $D=0
M1090 298 701 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=126860 $D=0
M1091 299 702 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=131490 $D=0
M1092 296 36 298 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=126860 $D=0
M1093 297 36 299 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=131490 $D=0
M1094 298 294 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=126860 $D=0
M1095 299 295 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=131490 $D=0
M1096 230 300 298 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=126860 $D=0
M1097 231 301 299 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=131490 $D=0
M1098 300 38 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=126860 $D=0
M1099 301 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=131490 $D=0
M1100 161 39 302 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=126860 $D=0
M1101 162 39 303 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=131490 $D=0
M1102 304 40 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=126860 $D=0
M1103 305 40 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=131490 $D=0
M1104 306 302 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=126860 $D=0
M1105 307 303 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=131490 $D=0
M1106 161 306 703 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=126860 $D=0
M1107 162 307 704 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=131490 $D=0
M1108 308 703 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=126860 $D=0
M1109 309 704 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=131490 $D=0
M1110 306 39 308 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=126860 $D=0
M1111 307 39 309 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=131490 $D=0
M1112 308 304 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=126860 $D=0
M1113 309 305 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=131490 $D=0
M1114 230 310 308 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=126860 $D=0
M1115 231 311 309 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=131490 $D=0
M1116 310 41 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=126860 $D=0
M1117 311 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=131490 $D=0
M1118 161 42 312 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=126860 $D=0
M1119 162 42 313 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=131490 $D=0
M1120 314 43 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=126860 $D=0
M1121 315 43 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=131490 $D=0
M1122 316 312 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=126860 $D=0
M1123 317 313 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=131490 $D=0
M1124 161 316 705 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=126860 $D=0
M1125 162 317 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=131490 $D=0
M1126 318 705 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=126860 $D=0
M1127 319 706 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=131490 $D=0
M1128 316 42 318 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=126860 $D=0
M1129 317 42 319 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=131490 $D=0
M1130 318 314 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=126860 $D=0
M1131 319 315 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=131490 $D=0
M1132 230 320 318 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=126860 $D=0
M1133 231 321 319 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=131490 $D=0
M1134 320 44 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=126860 $D=0
M1135 321 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=131490 $D=0
M1136 161 45 322 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=126860 $D=0
M1137 162 45 323 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=131490 $D=0
M1138 324 46 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=126860 $D=0
M1139 325 46 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=131490 $D=0
M1140 326 322 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=126860 $D=0
M1141 327 323 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=131490 $D=0
M1142 161 326 707 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=126860 $D=0
M1143 162 327 708 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=131490 $D=0
M1144 328 707 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=126860 $D=0
M1145 329 708 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=131490 $D=0
M1146 326 45 328 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=126860 $D=0
M1147 327 45 329 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=131490 $D=0
M1148 328 324 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=126860 $D=0
M1149 329 325 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=131490 $D=0
M1150 230 330 328 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=126860 $D=0
M1151 231 331 329 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=131490 $D=0
M1152 330 47 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=126860 $D=0
M1153 331 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=131490 $D=0
M1154 161 48 332 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=126860 $D=0
M1155 162 48 333 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=131490 $D=0
M1156 334 49 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=126860 $D=0
M1157 335 49 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=131490 $D=0
M1158 336 332 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=126860 $D=0
M1159 337 333 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=131490 $D=0
M1160 161 336 709 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=126860 $D=0
M1161 162 337 710 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=131490 $D=0
M1162 338 709 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=126860 $D=0
M1163 339 710 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=131490 $D=0
M1164 336 48 338 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=126860 $D=0
M1165 337 48 339 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=131490 $D=0
M1166 338 334 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=126860 $D=0
M1167 339 335 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=131490 $D=0
M1168 230 340 338 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=126860 $D=0
M1169 231 341 339 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=131490 $D=0
M1170 340 50 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=126860 $D=0
M1171 341 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=131490 $D=0
M1172 161 51 342 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=126860 $D=0
M1173 162 51 343 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=131490 $D=0
M1174 344 52 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=126860 $D=0
M1175 345 52 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=131490 $D=0
M1176 346 342 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=126860 $D=0
M1177 347 343 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=131490 $D=0
M1178 161 346 711 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=126860 $D=0
M1179 162 347 712 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=131490 $D=0
M1180 348 711 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=126860 $D=0
M1181 349 712 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=131490 $D=0
M1182 346 51 348 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=126860 $D=0
M1183 347 51 349 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=131490 $D=0
M1184 348 344 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=126860 $D=0
M1185 349 345 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=131490 $D=0
M1186 230 350 348 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=126860 $D=0
M1187 231 351 349 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=131490 $D=0
M1188 350 53 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=126860 $D=0
M1189 351 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=131490 $D=0
M1190 161 54 352 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=126860 $D=0
M1191 162 54 353 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=131490 $D=0
M1192 354 55 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=126860 $D=0
M1193 355 55 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=131490 $D=0
M1194 356 352 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=126860 $D=0
M1195 357 353 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=131490 $D=0
M1196 161 356 713 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=126860 $D=0
M1197 162 357 714 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=131490 $D=0
M1198 358 713 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=126860 $D=0
M1199 359 714 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=131490 $D=0
M1200 356 54 358 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=126860 $D=0
M1201 357 54 359 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=131490 $D=0
M1202 358 354 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=126860 $D=0
M1203 359 355 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=131490 $D=0
M1204 230 360 358 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=126860 $D=0
M1205 231 361 359 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=131490 $D=0
M1206 360 56 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=126860 $D=0
M1207 361 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=131490 $D=0
M1208 161 57 362 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=126860 $D=0
M1209 162 57 363 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=131490 $D=0
M1210 364 58 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=126860 $D=0
M1211 365 58 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=131490 $D=0
M1212 366 362 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=126860 $D=0
M1213 367 363 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=131490 $D=0
M1214 161 366 715 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=126860 $D=0
M1215 162 367 716 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=131490 $D=0
M1216 368 715 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=126860 $D=0
M1217 369 716 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=131490 $D=0
M1218 366 57 368 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=126860 $D=0
M1219 367 57 369 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=131490 $D=0
M1220 368 364 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=126860 $D=0
M1221 369 365 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=131490 $D=0
M1222 230 370 368 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=126860 $D=0
M1223 231 371 369 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=131490 $D=0
M1224 370 59 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=126860 $D=0
M1225 371 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=131490 $D=0
M1226 161 60 372 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=126860 $D=0
M1227 162 60 373 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=131490 $D=0
M1228 374 61 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=126860 $D=0
M1229 375 61 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=131490 $D=0
M1230 376 372 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=126860 $D=0
M1231 377 373 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=131490 $D=0
M1232 161 376 717 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=126860 $D=0
M1233 162 377 718 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=131490 $D=0
M1234 378 717 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=126860 $D=0
M1235 379 718 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=131490 $D=0
M1236 376 60 378 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=126860 $D=0
M1237 377 60 379 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=131490 $D=0
M1238 378 374 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=126860 $D=0
M1239 379 375 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=131490 $D=0
M1240 230 380 378 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=126860 $D=0
M1241 231 381 379 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=131490 $D=0
M1242 380 62 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=126860 $D=0
M1243 381 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=131490 $D=0
M1244 161 63 382 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=126860 $D=0
M1245 162 63 383 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=131490 $D=0
M1246 384 64 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=126860 $D=0
M1247 385 64 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=131490 $D=0
M1248 386 382 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=126860 $D=0
M1249 387 383 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=131490 $D=0
M1250 161 386 719 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=126860 $D=0
M1251 162 387 720 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=131490 $D=0
M1252 388 719 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=126860 $D=0
M1253 389 720 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=131490 $D=0
M1254 386 63 388 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=126860 $D=0
M1255 387 63 389 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=131490 $D=0
M1256 388 384 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=126860 $D=0
M1257 389 385 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=131490 $D=0
M1258 230 390 388 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=126860 $D=0
M1259 231 391 389 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=131490 $D=0
M1260 390 65 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=126860 $D=0
M1261 391 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=131490 $D=0
M1262 161 66 392 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=126860 $D=0
M1263 162 66 393 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=131490 $D=0
M1264 394 67 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=126860 $D=0
M1265 395 67 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=131490 $D=0
M1266 396 392 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=126860 $D=0
M1267 397 393 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=131490 $D=0
M1268 161 396 721 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=126860 $D=0
M1269 162 397 722 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=131490 $D=0
M1270 398 721 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=126860 $D=0
M1271 399 722 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=131490 $D=0
M1272 396 66 398 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=126860 $D=0
M1273 397 66 399 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=131490 $D=0
M1274 398 394 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=126860 $D=0
M1275 399 395 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=131490 $D=0
M1276 230 400 398 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=126860 $D=0
M1277 231 401 399 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=131490 $D=0
M1278 400 68 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=126860 $D=0
M1279 401 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=131490 $D=0
M1280 161 69 402 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=126860 $D=0
M1281 162 69 403 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=131490 $D=0
M1282 404 70 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=126860 $D=0
M1283 405 70 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=131490 $D=0
M1284 406 402 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=126860 $D=0
M1285 407 403 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=131490 $D=0
M1286 161 406 723 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=126860 $D=0
M1287 162 407 724 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=131490 $D=0
M1288 408 723 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=126860 $D=0
M1289 409 724 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=131490 $D=0
M1290 406 69 408 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=126860 $D=0
M1291 407 69 409 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=131490 $D=0
M1292 408 404 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=126860 $D=0
M1293 409 405 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=131490 $D=0
M1294 230 410 408 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=126860 $D=0
M1295 231 411 409 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=131490 $D=0
M1296 410 71 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=126860 $D=0
M1297 411 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=131490 $D=0
M1298 161 72 412 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=126860 $D=0
M1299 162 72 413 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=131490 $D=0
M1300 414 73 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=126860 $D=0
M1301 415 73 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=131490 $D=0
M1302 416 412 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=126860 $D=0
M1303 417 413 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=131490 $D=0
M1304 161 416 725 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=126860 $D=0
M1305 162 417 726 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=131490 $D=0
M1306 418 725 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=126860 $D=0
M1307 419 726 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=131490 $D=0
M1308 416 72 418 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=126860 $D=0
M1309 417 72 419 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=131490 $D=0
M1310 418 414 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=126860 $D=0
M1311 419 415 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=131490 $D=0
M1312 230 420 418 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=126860 $D=0
M1313 231 421 419 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=131490 $D=0
M1314 420 74 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=126860 $D=0
M1315 421 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=131490 $D=0
M1316 161 75 422 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=126860 $D=0
M1317 162 75 423 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=131490 $D=0
M1318 424 76 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=126860 $D=0
M1319 425 76 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=131490 $D=0
M1320 426 422 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=126860 $D=0
M1321 427 423 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=131490 $D=0
M1322 161 426 727 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=126860 $D=0
M1323 162 427 728 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=131490 $D=0
M1324 428 727 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=126860 $D=0
M1325 429 728 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=131490 $D=0
M1326 426 75 428 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=126860 $D=0
M1327 427 75 429 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=131490 $D=0
M1328 428 424 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=126860 $D=0
M1329 429 425 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=131490 $D=0
M1330 230 430 428 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=126860 $D=0
M1331 231 431 429 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=131490 $D=0
M1332 430 77 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=126860 $D=0
M1333 431 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=131490 $D=0
M1334 161 78 432 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=126860 $D=0
M1335 162 78 433 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=131490 $D=0
M1336 434 79 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=126860 $D=0
M1337 435 79 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=131490 $D=0
M1338 436 432 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=126860 $D=0
M1339 437 433 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=131490 $D=0
M1340 161 436 729 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=126860 $D=0
M1341 162 437 730 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=131490 $D=0
M1342 438 729 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=126860 $D=0
M1343 439 730 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=131490 $D=0
M1344 436 78 438 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=126860 $D=0
M1345 437 78 439 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=131490 $D=0
M1346 438 434 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=126860 $D=0
M1347 439 435 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=131490 $D=0
M1348 230 440 438 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=126860 $D=0
M1349 231 441 439 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=131490 $D=0
M1350 440 80 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=126860 $D=0
M1351 441 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=131490 $D=0
M1352 161 81 442 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=126860 $D=0
M1353 162 81 443 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=131490 $D=0
M1354 444 82 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=126860 $D=0
M1355 445 82 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=131490 $D=0
M1356 446 442 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=126860 $D=0
M1357 447 443 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=131490 $D=0
M1358 161 446 731 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=126860 $D=0
M1359 162 447 732 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=131490 $D=0
M1360 448 731 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=126860 $D=0
M1361 449 732 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=131490 $D=0
M1362 446 81 448 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=126860 $D=0
M1363 447 81 449 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=131490 $D=0
M1364 448 444 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=126860 $D=0
M1365 449 445 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=131490 $D=0
M1366 230 450 448 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=126860 $D=0
M1367 231 451 449 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=131490 $D=0
M1368 450 83 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=126860 $D=0
M1369 451 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=131490 $D=0
M1370 161 84 452 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=126860 $D=0
M1371 162 84 453 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=131490 $D=0
M1372 454 85 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=126860 $D=0
M1373 455 85 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=131490 $D=0
M1374 456 452 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=126860 $D=0
M1375 457 453 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=131490 $D=0
M1376 161 456 733 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=126860 $D=0
M1377 162 457 734 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=131490 $D=0
M1378 458 733 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=126860 $D=0
M1379 459 734 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=131490 $D=0
M1380 456 84 458 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=126860 $D=0
M1381 457 84 459 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=131490 $D=0
M1382 458 454 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=126860 $D=0
M1383 459 455 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=131490 $D=0
M1384 230 460 458 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=126860 $D=0
M1385 231 461 459 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=131490 $D=0
M1386 460 86 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=126860 $D=0
M1387 461 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=131490 $D=0
M1388 161 87 462 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=126860 $D=0
M1389 162 87 463 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=131490 $D=0
M1390 464 88 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=126860 $D=0
M1391 465 88 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=131490 $D=0
M1392 466 462 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=126860 $D=0
M1393 467 463 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=131490 $D=0
M1394 161 466 735 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=126860 $D=0
M1395 162 467 736 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=131490 $D=0
M1396 468 735 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=126860 $D=0
M1397 469 736 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=131490 $D=0
M1398 466 87 468 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=126860 $D=0
M1399 467 87 469 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=131490 $D=0
M1400 468 464 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=126860 $D=0
M1401 469 465 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=131490 $D=0
M1402 230 470 468 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=126860 $D=0
M1403 231 471 469 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=131490 $D=0
M1404 470 89 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=126860 $D=0
M1405 471 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=131490 $D=0
M1406 161 90 472 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=126860 $D=0
M1407 162 90 473 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=131490 $D=0
M1408 474 91 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=126860 $D=0
M1409 475 91 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=131490 $D=0
M1410 476 472 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=126860 $D=0
M1411 477 473 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=131490 $D=0
M1412 161 476 737 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=126860 $D=0
M1413 162 477 738 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=131490 $D=0
M1414 478 737 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=126860 $D=0
M1415 479 738 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=131490 $D=0
M1416 476 90 478 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=126860 $D=0
M1417 477 90 479 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=131490 $D=0
M1418 478 474 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=126860 $D=0
M1419 479 475 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=131490 $D=0
M1420 230 480 478 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=126860 $D=0
M1421 231 481 479 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=131490 $D=0
M1422 480 92 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=126860 $D=0
M1423 481 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=131490 $D=0
M1424 161 93 482 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=126860 $D=0
M1425 162 93 483 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=131490 $D=0
M1426 484 94 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=126860 $D=0
M1427 485 94 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=131490 $D=0
M1428 486 482 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=126860 $D=0
M1429 487 483 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=131490 $D=0
M1430 161 486 739 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=126860 $D=0
M1431 162 487 740 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=131490 $D=0
M1432 488 739 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=126860 $D=0
M1433 489 740 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=131490 $D=0
M1434 486 93 488 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=126860 $D=0
M1435 487 93 489 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=131490 $D=0
M1436 488 484 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=126860 $D=0
M1437 489 485 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=131490 $D=0
M1438 230 490 488 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=126860 $D=0
M1439 231 491 489 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=131490 $D=0
M1440 490 95 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=126860 $D=0
M1441 491 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=131490 $D=0
M1442 161 96 492 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=126860 $D=0
M1443 162 96 493 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=131490 $D=0
M1444 494 97 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=126860 $D=0
M1445 495 97 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=131490 $D=0
M1446 496 492 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=126860 $D=0
M1447 497 493 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=131490 $D=0
M1448 161 496 741 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=126860 $D=0
M1449 162 497 742 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=131490 $D=0
M1450 498 741 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=126860 $D=0
M1451 499 742 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=131490 $D=0
M1452 496 96 498 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=126860 $D=0
M1453 497 96 499 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=131490 $D=0
M1454 498 494 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=126860 $D=0
M1455 499 495 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=131490 $D=0
M1456 230 500 498 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=126860 $D=0
M1457 231 501 499 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=131490 $D=0
M1458 500 98 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=126860 $D=0
M1459 501 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=131490 $D=0
M1460 161 99 502 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=126860 $D=0
M1461 162 99 503 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=131490 $D=0
M1462 504 100 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=126860 $D=0
M1463 505 100 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=131490 $D=0
M1464 506 502 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=126860 $D=0
M1465 507 503 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=131490 $D=0
M1466 161 506 743 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=126860 $D=0
M1467 162 507 744 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=131490 $D=0
M1468 508 743 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=126860 $D=0
M1469 509 744 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=131490 $D=0
M1470 506 99 508 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=126860 $D=0
M1471 507 99 509 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=131490 $D=0
M1472 508 504 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=126860 $D=0
M1473 509 505 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=131490 $D=0
M1474 230 510 508 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=126860 $D=0
M1475 231 511 509 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=131490 $D=0
M1476 510 101 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=126860 $D=0
M1477 511 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=131490 $D=0
M1478 161 102 512 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=126860 $D=0
M1479 162 102 513 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=131490 $D=0
M1480 514 103 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=126860 $D=0
M1481 515 103 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=131490 $D=0
M1482 516 512 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=126860 $D=0
M1483 517 513 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=131490 $D=0
M1484 161 516 745 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=126860 $D=0
M1485 162 517 746 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=131490 $D=0
M1486 518 745 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=126860 $D=0
M1487 519 746 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=131490 $D=0
M1488 516 102 518 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=126860 $D=0
M1489 517 102 519 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=131490 $D=0
M1490 518 514 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=126860 $D=0
M1491 519 515 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=131490 $D=0
M1492 230 520 518 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=126860 $D=0
M1493 231 521 519 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=131490 $D=0
M1494 520 104 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=126860 $D=0
M1495 521 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=131490 $D=0
M1496 161 105 522 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=126860 $D=0
M1497 162 105 523 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=131490 $D=0
M1498 524 106 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=126860 $D=0
M1499 525 106 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=131490 $D=0
M1500 526 522 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=126860 $D=0
M1501 527 523 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=131490 $D=0
M1502 161 526 747 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=126860 $D=0
M1503 162 527 748 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=131490 $D=0
M1504 528 747 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=126860 $D=0
M1505 529 748 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=131490 $D=0
M1506 526 105 528 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=126860 $D=0
M1507 527 105 529 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=131490 $D=0
M1508 528 524 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=126860 $D=0
M1509 529 525 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=131490 $D=0
M1510 230 530 528 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=126860 $D=0
M1511 231 531 529 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=131490 $D=0
M1512 530 107 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=126860 $D=0
M1513 531 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=131490 $D=0
M1514 161 108 532 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=126860 $D=0
M1515 162 108 533 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=131490 $D=0
M1516 534 109 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=126860 $D=0
M1517 535 109 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=131490 $D=0
M1518 7 534 226 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=126860 $D=0
M1519 8 535 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=131490 $D=0
M1520 230 532 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=126860 $D=0
M1521 231 533 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=131490 $D=0
M1522 161 538 536 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=126860 $D=0
M1523 162 539 537 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=131490 $D=0
M1524 538 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=126860 $D=0
M1525 539 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=131490 $D=0
M1526 749 226 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=126860 $D=0
M1527 750 227 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=131490 $D=0
M1528 540 538 749 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=126860 $D=0
M1529 541 539 750 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=131490 $D=0
M1530 161 540 542 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=126860 $D=0
M1531 162 541 543 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=131490 $D=0
M1532 751 542 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=126860 $D=0
M1533 752 543 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=131490 $D=0
M1534 540 536 751 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=126860 $D=0
M1535 541 537 752 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=131490 $D=0
M1536 161 546 544 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=126860 $D=0
M1537 162 547 545 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=131490 $D=0
M1538 546 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=126860 $D=0
M1539 547 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=131490 $D=0
M1540 753 230 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=126860 $D=0
M1541 754 231 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=131490 $D=0
M1542 548 546 753 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=126860 $D=0
M1543 549 547 754 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=131490 $D=0
M1544 161 548 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=126860 $D=0
M1545 162 549 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=131490 $D=0
M1546 755 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=126860 $D=0
M1547 756 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=131490 $D=0
M1548 548 544 755 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=126860 $D=0
M1549 549 545 756 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=131490 $D=0
M1550 550 113 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=126860 $D=0
M1551 551 113 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=131490 $D=0
M1552 552 113 542 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=126860 $D=0
M1553 553 113 543 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=131490 $D=0
M1554 114 550 552 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=126860 $D=0
M1555 115 551 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=131490 $D=0
M1556 554 116 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=126860 $D=0
M1557 555 116 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=131490 $D=0
M1558 556 116 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=126860 $D=0
M1559 557 116 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=131490 $D=0
M1560 757 554 556 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=126860 $D=0
M1561 758 555 557 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=131490 $D=0
M1562 161 111 757 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=126860 $D=0
M1563 162 112 758 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=131490 $D=0
M1564 558 117 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=126860 $D=0
M1565 559 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=131490 $D=0
M1566 118 117 556 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=126860 $D=0
M1567 119 117 557 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=131490 $D=0
M1568 9 558 118 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=126860 $D=0
M1569 10 559 119 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=131490 $D=0
M1570 561 560 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=126860 $D=0
M1571 562 120 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=131490 $D=0
M1572 161 565 563 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=126860 $D=0
M1573 162 566 564 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=131490 $D=0
M1574 567 552 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=126860 $D=0
M1575 568 553 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=131490 $D=0
M1576 565 552 560 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=126860 $D=0
M1577 566 553 120 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=131490 $D=0
M1578 561 567 565 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=126860 $D=0
M1579 562 568 566 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=131490 $D=0
M1580 569 563 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=126860 $D=0
M1581 570 564 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=131490 $D=0
M1582 571 563 118 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=126860 $D=0
M1583 560 564 119 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=131490 $D=0
M1584 552 569 571 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=126860 $D=0
M1585 553 570 560 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=131490 $D=0
M1586 572 571 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=126860 $D=0
M1587 573 560 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=131490 $D=0
M1588 574 563 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=126860 $D=0
M1589 575 564 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=131490 $D=0
M1590 576 563 572 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=126860 $D=0
M1591 577 564 573 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=131490 $D=0
M1592 118 574 576 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=126860 $D=0
M1593 119 575 577 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=131490 $D=0
M1594 769 552 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=126500 $D=0
M1595 770 553 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=131130 $D=0
M1596 578 118 769 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=126500 $D=0
M1597 579 119 770 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=131130 $D=0
M1598 580 576 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=126860 $D=0
M1599 581 577 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=131490 $D=0
M1600 582 552 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=126860 $D=0
M1601 583 553 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=131490 $D=0
M1602 161 118 582 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=126860 $D=0
M1603 162 119 583 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=131490 $D=0
M1604 584 552 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=126860 $D=0
M1605 585 553 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=131490 $D=0
M1606 161 118 584 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=126860 $D=0
M1607 162 119 585 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=131490 $D=0
M1608 771 552 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=126680 $D=0
M1609 772 553 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=131310 $D=0
M1610 588 118 771 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=126680 $D=0
M1611 589 119 772 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=131310 $D=0
M1612 161 584 588 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=126860 $D=0
M1613 162 585 589 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=131490 $D=0
M1614 590 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=126860 $D=0
M1615 591 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=131490 $D=0
M1616 592 126 578 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=126860 $D=0
M1617 593 126 579 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=131490 $D=0
M1618 582 590 592 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=126860 $D=0
M1619 583 591 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=131490 $D=0
M1620 594 126 580 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=126860 $D=0
M1621 595 126 581 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=131490 $D=0
M1622 588 590 594 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=126860 $D=0
M1623 589 591 595 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=131490 $D=0
M1624 596 127 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=126860 $D=0
M1625 597 127 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=131490 $D=0
M1626 598 127 594 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=126860 $D=0
M1627 599 127 595 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=131490 $D=0
M1628 592 596 598 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=126860 $D=0
M1629 593 597 599 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=131490 $D=0
M1630 11 598 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=126860 $D=0
M1631 12 599 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=131490 $D=0
M1632 600 129 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=126860 $D=0
M1633 601 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=131490 $D=0
M1634 602 129 130 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=126860 $D=0
M1635 603 129 131 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=131490 $D=0
M1636 132 600 602 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=126860 $D=0
M1637 133 601 603 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=131490 $D=0
M1638 604 129 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=126860 $D=0
M1639 605 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=131490 $D=0
M1640 606 129 134 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=126860 $D=0
M1641 607 129 135 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=131490 $D=0
M1642 136 604 606 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=126860 $D=0
M1643 137 605 607 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=131490 $D=0
M1644 608 129 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=126860 $D=0
M1645 609 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=131490 $D=0
M1646 138 129 123 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=126860 $D=0
M1647 138 129 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=131490 $D=0
M1648 128 608 138 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=126860 $D=0
M1649 139 609 138 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=131490 $D=0
M1650 610 129 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=126860 $D=0
M1651 611 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=131490 $D=0
M1652 612 129 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=126860 $D=0
M1653 613 129 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=131490 $D=0
M1654 140 610 612 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=126860 $D=0
M1655 141 611 613 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=131490 $D=0
M1656 614 129 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=126860 $D=0
M1657 615 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=131490 $D=0
M1658 616 129 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=126860 $D=0
M1659 617 129 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=131490 $D=0
M1660 142 614 616 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=126860 $D=0
M1661 143 615 617 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=131490 $D=0
M1662 161 552 759 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=126860 $D=0
M1663 162 553 760 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=131490 $D=0
M1664 133 759 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=126860 $D=0
M1665 130 760 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=131490 $D=0
M1666 618 144 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=126860 $D=0
M1667 619 144 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=131490 $D=0
M1668 145 144 133 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=126860 $D=0
M1669 146 144 130 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=131490 $D=0
M1670 602 618 145 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=126860 $D=0
M1671 603 619 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=131490 $D=0
M1672 620 147 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=126860 $D=0
M1673 621 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=131490 $D=0
M1674 148 147 145 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=126860 $D=0
M1675 125 147 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=131490 $D=0
M1676 606 620 148 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=126860 $D=0
M1677 607 621 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=131490 $D=0
M1678 622 149 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=126860 $D=0
M1679 623 149 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=131490 $D=0
M1680 121 149 148 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=126860 $D=0
M1681 122 149 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=131490 $D=0
M1682 138 622 121 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=126860 $D=0
M1683 138 623 122 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=131490 $D=0
M1684 624 119 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=126860 $D=0
M1685 625 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=131490 $D=0
M1686 150 119 121 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=126860 $D=0
M1687 151 119 122 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=131490 $D=0
M1688 612 624 150 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=126860 $D=0
M1689 613 625 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=131490 $D=0
M1690 626 118 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=126860 $D=0
M1691 627 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=131490 $D=0
M1692 202 118 150 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=126860 $D=0
M1693 203 118 151 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=131490 $D=0
M1694 616 626 202 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=126860 $D=0
M1695 617 627 203 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=131490 $D=0
M1696 628 152 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=126860 $D=0
M1697 629 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=131490 $D=0
M1698 630 152 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=126860 $D=0
M1699 631 152 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=131490 $D=0
M1700 9 628 630 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=126860 $D=0
M1701 10 629 631 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=131490 $D=0
M1702 632 542 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=126860 $D=0
M1703 633 543 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=131490 $D=0
M1704 161 630 632 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=126860 $D=0
M1705 162 631 633 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=131490 $D=0
M1706 773 542 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=126680 $D=0
M1707 774 543 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=131310 $D=0
M1708 636 630 773 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=126680 $D=0
M1709 637 631 774 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=131310 $D=0
M1710 161 632 636 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=126860 $D=0
M1711 162 633 637 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=131490 $D=0
M1712 761 153 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=126860 $D=0
M1713 762 638 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=131490 $D=0
M1714 161 636 761 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=126860 $D=0
M1715 162 637 762 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=131490 $D=0
M1716 638 761 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=126860 $D=0
M1717 154 762 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=131490 $D=0
M1718 775 542 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=126500 $D=0
M1719 776 543 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=131130 $D=0
M1720 639 641 775 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=126500 $D=0
M1721 640 642 776 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=131130 $D=0
M1722 641 630 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=126860 $D=0
M1723 642 631 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=131490 $D=0
M1724 643 639 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=126860 $D=0
M1725 644 640 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=131490 $D=0
M1726 161 153 643 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=126860 $D=0
M1727 162 638 644 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=131490 $D=0
M1728 646 155 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=126860 $D=0
M1729 647 645 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=131490 $D=0
M1730 645 643 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=126860 $D=0
M1731 156 644 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=131490 $D=0
M1732 161 646 645 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=126860 $D=0
M1733 162 647 156 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=131490 $D=0
M1734 649 648 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=126860 $D=0
M1735 650 157 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=131490 $D=0
M1736 161 653 651 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=126860 $D=0
M1737 162 654 652 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=131490 $D=0
M1738 655 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=126860 $D=0
M1739 656 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=131490 $D=0
M1740 653 114 648 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=126860 $D=0
M1741 654 115 157 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=131490 $D=0
M1742 649 655 653 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=126860 $D=0
M1743 650 656 654 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=131490 $D=0
M1744 657 651 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=126860 $D=0
M1745 658 652 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=131490 $D=0
M1746 158 651 7 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=126860 $D=0
M1747 648 652 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=131490 $D=0
M1748 114 657 158 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=126860 $D=0
M1749 115 658 648 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=131490 $D=0
M1750 659 158 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=126860 $D=0
M1751 660 648 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=131490 $D=0
M1752 661 651 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=126860 $D=0
M1753 662 652 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=131490 $D=0
M1754 204 651 659 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=126860 $D=0
M1755 205 652 660 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=131490 $D=0
M1756 7 661 204 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=126860 $D=0
M1757 8 662 205 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=131490 $D=0
M1758 663 159 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=126860 $D=0
M1759 664 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=131490 $D=0
M1760 665 159 204 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=126860 $D=0
M1761 666 159 205 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=131490 $D=0
M1762 11 663 665 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=126860 $D=0
M1763 12 664 666 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=131490 $D=0
M1764 667 160 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=126860 $D=0
M1765 668 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=131490 $D=0
M1766 160 160 665 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=126860 $D=0
M1767 160 160 666 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=131490 $D=0
M1768 7 667 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=126860 $D=0
M1769 8 668 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=131490 $D=0
M1770 669 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=126860 $D=0
M1771 670 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=131490 $D=0
M1772 161 669 671 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=126860 $D=0
M1773 162 670 672 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=131490 $D=0
M1774 673 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=126860 $D=0
M1775 674 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=131490 $D=0
M1776 675 671 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=126860 $D=0
M1777 676 672 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=131490 $D=0
M1778 161 675 763 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=126860 $D=0
M1779 162 676 764 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=131490 $D=0
M1780 677 763 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=126860 $D=0
M1781 678 764 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=131490 $D=0
M1782 675 669 677 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=126860 $D=0
M1783 676 670 678 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=131490 $D=0
M1784 679 673 677 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=126860 $D=0
M1785 680 674 678 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=131490 $D=0
M1786 161 683 681 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=126860 $D=0
M1787 162 684 682 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=131490 $D=0
M1788 683 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=126860 $D=0
M1789 684 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=131490 $D=0
M1790 765 679 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=126860 $D=0
M1791 766 680 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=131490 $D=0
M1792 685 683 765 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=126860 $D=0
M1793 686 684 766 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=131490 $D=0
M1794 161 685 114 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=126860 $D=0
M1795 162 686 115 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=131490 $D=0
M1796 767 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=126860 $D=0
M1797 768 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=131490 $D=0
M1798 685 681 767 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=126860 $D=0
M1799 686 682 768 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=131490 $D=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164
** N=799 EP=163 IP=1514 FDC=1800
M0 188 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=116350 $D=1
M1 189 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=120980 $D=1
M2 190 188 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=116350 $D=1
M3 191 189 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=120980 $D=1
M4 7 1 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=116350 $D=1
M5 8 1 191 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=120980 $D=1
M6 192 188 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=116350 $D=1
M7 193 189 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=120980 $D=1
M8 2 1 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=116350 $D=1
M9 3 1 193 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=120980 $D=1
M10 194 188 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=116350 $D=1
M11 195 189 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=120980 $D=1
M12 2 1 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=116350 $D=1
M13 3 1 195 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=120980 $D=1
M14 198 196 194 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=116350 $D=1
M15 199 197 195 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=120980 $D=1
M16 196 4 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=116350 $D=1
M17 197 4 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=120980 $D=1
M18 200 196 192 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=116350 $D=1
M19 201 197 193 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=120980 $D=1
M20 190 4 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=116350 $D=1
M21 191 4 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=120980 $D=1
M22 202 5 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=116350 $D=1
M23 203 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=120980 $D=1
M24 204 202 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=116350 $D=1
M25 205 203 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=120980 $D=1
M26 198 5 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=116350 $D=1
M27 199 5 205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=120980 $D=1
M28 206 6 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=116350 $D=1
M29 207 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=120980 $D=1
M30 208 206 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=116350 $D=1
M31 209 207 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=120980 $D=1
M32 9 6 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=116350 $D=1
M33 10 6 209 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=120980 $D=1
M34 210 206 11 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=116350 $D=1
M35 211 207 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=120980 $D=1
M36 212 6 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=116350 $D=1
M37 213 6 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=120980 $D=1
M38 216 206 214 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=116350 $D=1
M39 217 207 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=120980 $D=1
M40 204 6 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=116350 $D=1
M41 205 6 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=120980 $D=1
M42 220 218 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=116350 $D=1
M43 221 219 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=120980 $D=1
M44 218 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=116350 $D=1
M45 219 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=120980 $D=1
M46 222 218 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=116350 $D=1
M47 223 219 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=120980 $D=1
M48 208 13 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=116350 $D=1
M49 209 13 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=120980 $D=1
M50 224 14 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=116350 $D=1
M51 225 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=120980 $D=1
M52 226 224 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=116350 $D=1
M53 227 225 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=120980 $D=1
M54 220 14 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=116350 $D=1
M55 221 14 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=120980 $D=1
M56 7 15 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=116350 $D=1
M57 8 15 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=120980 $D=1
M58 230 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=116350 $D=1
M59 231 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=120980 $D=1
M60 232 15 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=116350 $D=1
M61 233 15 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=120980 $D=1
M62 7 232 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=116350 $D=1
M63 8 233 699 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=120980 $D=1
M64 234 698 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=116350 $D=1
M65 235 699 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=120980 $D=1
M66 232 228 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=116350 $D=1
M67 233 229 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=120980 $D=1
M68 234 16 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=116350 $D=1
M69 235 16 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=120980 $D=1
M70 240 17 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=116350 $D=1
M71 241 17 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=120980 $D=1
M72 238 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=116350 $D=1
M73 239 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=120980 $D=1
M74 7 18 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=116350 $D=1
M75 8 18 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=120980 $D=1
M76 244 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=116350 $D=1
M77 245 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=120980 $D=1
M78 246 18 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=116350 $D=1
M79 247 18 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=120980 $D=1
M80 7 246 700 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=116350 $D=1
M81 8 247 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=120980 $D=1
M82 248 700 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=116350 $D=1
M83 249 701 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=120980 $D=1
M84 246 242 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=116350 $D=1
M85 247 243 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=120980 $D=1
M86 248 19 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=116350 $D=1
M87 249 19 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=120980 $D=1
M88 240 20 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=116350 $D=1
M89 241 20 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=120980 $D=1
M90 250 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=116350 $D=1
M91 251 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=120980 $D=1
M92 7 21 252 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=116350 $D=1
M93 8 21 253 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=120980 $D=1
M94 254 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=116350 $D=1
M95 255 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=120980 $D=1
M96 256 21 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=116350 $D=1
M97 257 21 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=120980 $D=1
M98 7 256 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=116350 $D=1
M99 8 257 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=120980 $D=1
M100 258 702 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=116350 $D=1
M101 259 703 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=120980 $D=1
M102 256 252 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=116350 $D=1
M103 257 253 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=120980 $D=1
M104 258 22 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=116350 $D=1
M105 259 22 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=120980 $D=1
M106 240 23 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=116350 $D=1
M107 241 23 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=120980 $D=1
M108 260 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=116350 $D=1
M109 261 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=120980 $D=1
M110 7 24 262 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=116350 $D=1
M111 8 24 263 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=120980 $D=1
M112 264 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=116350 $D=1
M113 265 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=120980 $D=1
M114 266 24 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=116350 $D=1
M115 267 24 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=120980 $D=1
M116 7 266 704 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=116350 $D=1
M117 8 267 705 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=120980 $D=1
M118 268 704 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=116350 $D=1
M119 269 705 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=120980 $D=1
M120 266 262 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=116350 $D=1
M121 267 263 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=120980 $D=1
M122 268 25 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=116350 $D=1
M123 269 25 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=120980 $D=1
M124 240 26 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=116350 $D=1
M125 241 26 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=120980 $D=1
M126 270 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=116350 $D=1
M127 271 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=120980 $D=1
M128 7 27 272 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=116350 $D=1
M129 8 27 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=120980 $D=1
M130 274 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=116350 $D=1
M131 275 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=120980 $D=1
M132 276 27 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=116350 $D=1
M133 277 27 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=120980 $D=1
M134 7 276 706 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=116350 $D=1
M135 8 277 707 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=120980 $D=1
M136 278 706 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=116350 $D=1
M137 279 707 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=120980 $D=1
M138 276 272 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=116350 $D=1
M139 277 273 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=120980 $D=1
M140 278 28 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=116350 $D=1
M141 279 28 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=120980 $D=1
M142 240 29 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=116350 $D=1
M143 241 29 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=120980 $D=1
M144 280 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=116350 $D=1
M145 281 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=120980 $D=1
M146 7 30 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=116350 $D=1
M147 8 30 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=120980 $D=1
M148 284 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=116350 $D=1
M149 285 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=120980 $D=1
M150 286 30 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=116350 $D=1
M151 287 30 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=120980 $D=1
M152 7 286 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=116350 $D=1
M153 8 287 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=120980 $D=1
M154 288 708 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=116350 $D=1
M155 289 709 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=120980 $D=1
M156 286 282 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=116350 $D=1
M157 287 283 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=120980 $D=1
M158 288 31 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=116350 $D=1
M159 289 31 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=120980 $D=1
M160 240 32 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=116350 $D=1
M161 241 32 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=120980 $D=1
M162 290 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=116350 $D=1
M163 291 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=120980 $D=1
M164 7 33 292 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=116350 $D=1
M165 8 33 293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=120980 $D=1
M166 294 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=116350 $D=1
M167 295 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=120980 $D=1
M168 296 33 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=116350 $D=1
M169 297 33 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=120980 $D=1
M170 7 296 710 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=116350 $D=1
M171 8 297 711 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=120980 $D=1
M172 298 710 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=116350 $D=1
M173 299 711 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=120980 $D=1
M174 296 292 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=116350 $D=1
M175 297 293 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=120980 $D=1
M176 298 34 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=116350 $D=1
M177 299 34 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=120980 $D=1
M178 240 35 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=116350 $D=1
M179 241 35 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=120980 $D=1
M180 300 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=116350 $D=1
M181 301 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=120980 $D=1
M182 7 36 302 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=116350 $D=1
M183 8 36 303 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=120980 $D=1
M184 304 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=116350 $D=1
M185 305 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=120980 $D=1
M186 306 36 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=116350 $D=1
M187 307 36 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=120980 $D=1
M188 7 306 712 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=116350 $D=1
M189 8 307 713 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=120980 $D=1
M190 308 712 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=116350 $D=1
M191 309 713 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=120980 $D=1
M192 306 302 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=116350 $D=1
M193 307 303 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=120980 $D=1
M194 308 37 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=116350 $D=1
M195 309 37 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=120980 $D=1
M196 240 38 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=116350 $D=1
M197 241 38 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=120980 $D=1
M198 310 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=116350 $D=1
M199 311 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=120980 $D=1
M200 7 39 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=116350 $D=1
M201 8 39 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=120980 $D=1
M202 314 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=116350 $D=1
M203 315 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=120980 $D=1
M204 316 39 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=116350 $D=1
M205 317 39 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=120980 $D=1
M206 7 316 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=116350 $D=1
M207 8 317 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=120980 $D=1
M208 318 714 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=116350 $D=1
M209 319 715 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=120980 $D=1
M210 316 312 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=116350 $D=1
M211 317 313 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=120980 $D=1
M212 318 40 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=116350 $D=1
M213 319 40 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=120980 $D=1
M214 240 41 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=116350 $D=1
M215 241 41 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=120980 $D=1
M216 320 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=116350 $D=1
M217 321 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=120980 $D=1
M218 7 42 322 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=116350 $D=1
M219 8 42 323 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=120980 $D=1
M220 324 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=116350 $D=1
M221 325 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=120980 $D=1
M222 326 42 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=116350 $D=1
M223 327 42 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=120980 $D=1
M224 7 326 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=116350 $D=1
M225 8 327 717 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=120980 $D=1
M226 328 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=116350 $D=1
M227 329 717 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=120980 $D=1
M228 326 322 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=116350 $D=1
M229 327 323 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=120980 $D=1
M230 328 43 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=116350 $D=1
M231 329 43 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=120980 $D=1
M232 240 44 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=116350 $D=1
M233 241 44 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=120980 $D=1
M234 330 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=116350 $D=1
M235 331 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=120980 $D=1
M236 7 45 332 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=116350 $D=1
M237 8 45 333 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=120980 $D=1
M238 334 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=116350 $D=1
M239 335 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=120980 $D=1
M240 336 45 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=116350 $D=1
M241 337 45 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=120980 $D=1
M242 7 336 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=116350 $D=1
M243 8 337 719 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=120980 $D=1
M244 338 718 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=116350 $D=1
M245 339 719 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=120980 $D=1
M246 336 332 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=116350 $D=1
M247 337 333 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=120980 $D=1
M248 338 46 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=116350 $D=1
M249 339 46 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=120980 $D=1
M250 240 47 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=116350 $D=1
M251 241 47 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=120980 $D=1
M252 340 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=116350 $D=1
M253 341 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=120980 $D=1
M254 7 48 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=116350 $D=1
M255 8 48 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=120980 $D=1
M256 344 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=116350 $D=1
M257 345 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=120980 $D=1
M258 346 48 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=116350 $D=1
M259 347 48 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=120980 $D=1
M260 7 346 720 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=116350 $D=1
M261 8 347 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=120980 $D=1
M262 348 720 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=116350 $D=1
M263 349 721 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=120980 $D=1
M264 346 342 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=116350 $D=1
M265 347 343 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=120980 $D=1
M266 348 49 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=116350 $D=1
M267 349 49 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=120980 $D=1
M268 240 50 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=116350 $D=1
M269 241 50 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=120980 $D=1
M270 350 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=116350 $D=1
M271 351 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=120980 $D=1
M272 7 51 352 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=116350 $D=1
M273 8 51 353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=120980 $D=1
M274 354 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=116350 $D=1
M275 355 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=120980 $D=1
M276 356 51 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=116350 $D=1
M277 357 51 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=120980 $D=1
M278 7 356 722 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=116350 $D=1
M279 8 357 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=120980 $D=1
M280 358 722 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=116350 $D=1
M281 359 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=120980 $D=1
M282 356 352 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=116350 $D=1
M283 357 353 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=120980 $D=1
M284 358 52 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=116350 $D=1
M285 359 52 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=120980 $D=1
M286 240 53 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=116350 $D=1
M287 241 53 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=120980 $D=1
M288 360 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=116350 $D=1
M289 361 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=120980 $D=1
M290 7 54 362 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=116350 $D=1
M291 8 54 363 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=120980 $D=1
M292 364 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=116350 $D=1
M293 365 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=120980 $D=1
M294 366 54 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=116350 $D=1
M295 367 54 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=120980 $D=1
M296 7 366 724 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=116350 $D=1
M297 8 367 725 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=120980 $D=1
M298 368 724 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=116350 $D=1
M299 369 725 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=120980 $D=1
M300 366 362 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=116350 $D=1
M301 367 363 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=120980 $D=1
M302 368 55 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=116350 $D=1
M303 369 55 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=120980 $D=1
M304 240 56 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=116350 $D=1
M305 241 56 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=120980 $D=1
M306 370 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=116350 $D=1
M307 371 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=120980 $D=1
M308 7 57 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=116350 $D=1
M309 8 57 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=120980 $D=1
M310 374 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=116350 $D=1
M311 375 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=120980 $D=1
M312 376 57 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=116350 $D=1
M313 377 57 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=120980 $D=1
M314 7 376 726 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=116350 $D=1
M315 8 377 727 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=120980 $D=1
M316 378 726 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=116350 $D=1
M317 379 727 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=120980 $D=1
M318 376 372 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=116350 $D=1
M319 377 373 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=120980 $D=1
M320 378 58 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=116350 $D=1
M321 379 58 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=120980 $D=1
M322 240 59 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=116350 $D=1
M323 241 59 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=120980 $D=1
M324 380 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=116350 $D=1
M325 381 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=120980 $D=1
M326 7 60 382 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=116350 $D=1
M327 8 60 383 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=120980 $D=1
M328 384 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=116350 $D=1
M329 385 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=120980 $D=1
M330 386 60 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=116350 $D=1
M331 387 60 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=120980 $D=1
M332 7 386 728 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=116350 $D=1
M333 8 387 729 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=120980 $D=1
M334 388 728 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=116350 $D=1
M335 389 729 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=120980 $D=1
M336 386 382 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=116350 $D=1
M337 387 383 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=120980 $D=1
M338 388 61 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=116350 $D=1
M339 389 61 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=120980 $D=1
M340 240 62 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=116350 $D=1
M341 241 62 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=120980 $D=1
M342 390 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=116350 $D=1
M343 391 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=120980 $D=1
M344 7 63 392 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=116350 $D=1
M345 8 63 393 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=120980 $D=1
M346 394 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=116350 $D=1
M347 395 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=120980 $D=1
M348 396 63 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=116350 $D=1
M349 397 63 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=120980 $D=1
M350 7 396 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=116350 $D=1
M351 8 397 731 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=120980 $D=1
M352 398 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=116350 $D=1
M353 399 731 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=120980 $D=1
M354 396 392 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=116350 $D=1
M355 397 393 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=120980 $D=1
M356 398 64 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=116350 $D=1
M357 399 64 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=120980 $D=1
M358 240 65 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=116350 $D=1
M359 241 65 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=120980 $D=1
M360 400 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=116350 $D=1
M361 401 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=120980 $D=1
M362 7 66 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=116350 $D=1
M363 8 66 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=120980 $D=1
M364 404 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=116350 $D=1
M365 405 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=120980 $D=1
M366 406 66 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=116350 $D=1
M367 407 66 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=120980 $D=1
M368 7 406 732 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=116350 $D=1
M369 8 407 733 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=120980 $D=1
M370 408 732 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=116350 $D=1
M371 409 733 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=120980 $D=1
M372 406 402 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=116350 $D=1
M373 407 403 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=120980 $D=1
M374 408 67 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=116350 $D=1
M375 409 67 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=120980 $D=1
M376 240 68 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=116350 $D=1
M377 241 68 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=120980 $D=1
M378 410 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=116350 $D=1
M379 411 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=120980 $D=1
M380 7 69 412 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=116350 $D=1
M381 8 69 413 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=120980 $D=1
M382 414 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=116350 $D=1
M383 415 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=120980 $D=1
M384 416 69 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=116350 $D=1
M385 417 69 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=120980 $D=1
M386 7 416 734 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=116350 $D=1
M387 8 417 735 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=120980 $D=1
M388 418 734 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=116350 $D=1
M389 419 735 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=120980 $D=1
M390 416 412 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=116350 $D=1
M391 417 413 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=120980 $D=1
M392 418 70 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=116350 $D=1
M393 419 70 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=120980 $D=1
M394 240 71 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=116350 $D=1
M395 241 71 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=120980 $D=1
M396 420 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=116350 $D=1
M397 421 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=120980 $D=1
M398 7 72 422 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=116350 $D=1
M399 8 72 423 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=120980 $D=1
M400 424 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=116350 $D=1
M401 425 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=120980 $D=1
M402 426 72 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=116350 $D=1
M403 427 72 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=120980 $D=1
M404 7 426 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=116350 $D=1
M405 8 427 737 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=120980 $D=1
M406 428 736 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=116350 $D=1
M407 429 737 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=120980 $D=1
M408 426 422 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=116350 $D=1
M409 427 423 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=120980 $D=1
M410 428 73 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=116350 $D=1
M411 429 73 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=120980 $D=1
M412 240 74 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=116350 $D=1
M413 241 74 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=120980 $D=1
M414 430 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=116350 $D=1
M415 431 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=120980 $D=1
M416 7 75 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=116350 $D=1
M417 8 75 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=120980 $D=1
M418 434 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=116350 $D=1
M419 435 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=120980 $D=1
M420 436 75 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=116350 $D=1
M421 437 75 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=120980 $D=1
M422 7 436 738 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=116350 $D=1
M423 8 437 739 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=120980 $D=1
M424 438 738 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=116350 $D=1
M425 439 739 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=120980 $D=1
M426 436 432 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=116350 $D=1
M427 437 433 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=120980 $D=1
M428 438 76 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=116350 $D=1
M429 439 76 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=120980 $D=1
M430 240 77 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=116350 $D=1
M431 241 77 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=120980 $D=1
M432 440 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=116350 $D=1
M433 441 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=120980 $D=1
M434 7 78 442 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=116350 $D=1
M435 8 78 443 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=120980 $D=1
M436 444 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=116350 $D=1
M437 445 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=120980 $D=1
M438 446 78 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=116350 $D=1
M439 447 78 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=120980 $D=1
M440 7 446 740 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=116350 $D=1
M441 8 447 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=120980 $D=1
M442 448 740 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=116350 $D=1
M443 449 741 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=120980 $D=1
M444 446 442 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=116350 $D=1
M445 447 443 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=120980 $D=1
M446 448 79 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=116350 $D=1
M447 449 79 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=120980 $D=1
M448 240 80 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=116350 $D=1
M449 241 80 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=120980 $D=1
M450 450 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=116350 $D=1
M451 451 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=120980 $D=1
M452 7 81 452 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=116350 $D=1
M453 8 81 453 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=120980 $D=1
M454 454 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=116350 $D=1
M455 455 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=120980 $D=1
M456 456 81 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=116350 $D=1
M457 457 81 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=120980 $D=1
M458 7 456 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=116350 $D=1
M459 8 457 743 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=120980 $D=1
M460 458 742 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=116350 $D=1
M461 459 743 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=120980 $D=1
M462 456 452 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=116350 $D=1
M463 457 453 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=120980 $D=1
M464 458 82 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=116350 $D=1
M465 459 82 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=120980 $D=1
M466 240 83 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=116350 $D=1
M467 241 83 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=120980 $D=1
M468 460 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=116350 $D=1
M469 461 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=120980 $D=1
M470 7 84 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=116350 $D=1
M471 8 84 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=120980 $D=1
M472 464 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=116350 $D=1
M473 465 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=120980 $D=1
M474 466 84 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=116350 $D=1
M475 467 84 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=120980 $D=1
M476 7 466 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=116350 $D=1
M477 8 467 745 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=120980 $D=1
M478 468 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=116350 $D=1
M479 469 745 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=120980 $D=1
M480 466 462 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=116350 $D=1
M481 467 463 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=120980 $D=1
M482 468 85 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=116350 $D=1
M483 469 85 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=120980 $D=1
M484 240 86 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=116350 $D=1
M485 241 86 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=120980 $D=1
M486 470 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=116350 $D=1
M487 471 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=120980 $D=1
M488 7 87 472 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=116350 $D=1
M489 8 87 473 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=120980 $D=1
M490 474 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=116350 $D=1
M491 475 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=120980 $D=1
M492 476 87 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=116350 $D=1
M493 477 87 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=120980 $D=1
M494 7 476 746 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=116350 $D=1
M495 8 477 747 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=120980 $D=1
M496 478 746 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=116350 $D=1
M497 479 747 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=120980 $D=1
M498 476 472 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=116350 $D=1
M499 477 473 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=120980 $D=1
M500 478 88 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=116350 $D=1
M501 479 88 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=120980 $D=1
M502 240 89 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=116350 $D=1
M503 241 89 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=120980 $D=1
M504 480 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=116350 $D=1
M505 481 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=120980 $D=1
M506 7 90 482 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=116350 $D=1
M507 8 90 483 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=120980 $D=1
M508 484 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=116350 $D=1
M509 485 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=120980 $D=1
M510 486 90 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=116350 $D=1
M511 487 90 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=120980 $D=1
M512 7 486 748 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=116350 $D=1
M513 8 487 749 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=120980 $D=1
M514 488 748 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=116350 $D=1
M515 489 749 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=120980 $D=1
M516 486 482 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=116350 $D=1
M517 487 483 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=120980 $D=1
M518 488 91 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=116350 $D=1
M519 489 91 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=120980 $D=1
M520 240 92 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=116350 $D=1
M521 241 92 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=120980 $D=1
M522 490 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=116350 $D=1
M523 491 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=120980 $D=1
M524 7 93 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=116350 $D=1
M525 8 93 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=120980 $D=1
M526 494 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=116350 $D=1
M527 495 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=120980 $D=1
M528 496 93 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=116350 $D=1
M529 497 93 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=120980 $D=1
M530 7 496 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=116350 $D=1
M531 8 497 751 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=120980 $D=1
M532 498 750 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=116350 $D=1
M533 499 751 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=120980 $D=1
M534 496 492 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=116350 $D=1
M535 497 493 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=120980 $D=1
M536 498 94 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=116350 $D=1
M537 499 94 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=120980 $D=1
M538 240 95 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=116350 $D=1
M539 241 95 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=120980 $D=1
M540 500 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=116350 $D=1
M541 501 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=120980 $D=1
M542 7 96 502 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=116350 $D=1
M543 8 96 503 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=120980 $D=1
M544 504 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=116350 $D=1
M545 505 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=120980 $D=1
M546 506 96 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=116350 $D=1
M547 507 96 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=120980 $D=1
M548 7 506 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=116350 $D=1
M549 8 507 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=120980 $D=1
M550 508 752 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=116350 $D=1
M551 509 753 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=120980 $D=1
M552 506 502 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=116350 $D=1
M553 507 503 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=120980 $D=1
M554 508 97 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=116350 $D=1
M555 509 97 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=120980 $D=1
M556 240 98 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=116350 $D=1
M557 241 98 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=120980 $D=1
M558 510 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=116350 $D=1
M559 511 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=120980 $D=1
M560 7 99 512 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=116350 $D=1
M561 8 99 513 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=120980 $D=1
M562 514 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=116350 $D=1
M563 515 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=120980 $D=1
M564 516 99 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=116350 $D=1
M565 517 99 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=120980 $D=1
M566 7 516 754 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=116350 $D=1
M567 8 517 755 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=120980 $D=1
M568 518 754 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=116350 $D=1
M569 519 755 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=120980 $D=1
M570 516 512 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=116350 $D=1
M571 517 513 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=120980 $D=1
M572 518 100 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=116350 $D=1
M573 519 100 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=120980 $D=1
M574 240 101 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=116350 $D=1
M575 241 101 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=120980 $D=1
M576 520 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=116350 $D=1
M577 521 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=120980 $D=1
M578 7 102 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=116350 $D=1
M579 8 102 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=120980 $D=1
M580 524 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=116350 $D=1
M581 525 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=120980 $D=1
M582 526 102 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=116350 $D=1
M583 527 102 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=120980 $D=1
M584 7 526 756 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=116350 $D=1
M585 8 527 757 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=120980 $D=1
M586 528 756 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=116350 $D=1
M587 529 757 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=120980 $D=1
M588 526 522 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=116350 $D=1
M589 527 523 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=120980 $D=1
M590 528 103 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=116350 $D=1
M591 529 103 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=120980 $D=1
M592 240 104 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=116350 $D=1
M593 241 104 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=120980 $D=1
M594 530 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=116350 $D=1
M595 531 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=120980 $D=1
M596 7 105 532 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=116350 $D=1
M597 8 105 533 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=120980 $D=1
M598 534 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=116350 $D=1
M599 535 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=120980 $D=1
M600 536 105 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=116350 $D=1
M601 537 105 227 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=120980 $D=1
M602 7 536 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=116350 $D=1
M603 8 537 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=120980 $D=1
M604 538 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=116350 $D=1
M605 539 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=120980 $D=1
M606 536 532 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=116350 $D=1
M607 537 533 539 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=120980 $D=1
M608 538 106 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=116350 $D=1
M609 539 106 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=120980 $D=1
M610 240 107 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=116350 $D=1
M611 241 107 539 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=120980 $D=1
M612 540 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=116350 $D=1
M613 541 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=120980 $D=1
M614 7 108 542 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=116350 $D=1
M615 8 108 543 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=120980 $D=1
M616 544 109 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=116350 $D=1
M617 545 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=120980 $D=1
M618 7 109 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=116350 $D=1
M619 8 109 237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=120980 $D=1
M620 240 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=116350 $D=1
M621 241 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=120980 $D=1
M622 7 548 546 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=116350 $D=1
M623 8 549 547 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=120980 $D=1
M624 548 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=116350 $D=1
M625 549 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=120980 $D=1
M626 760 236 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=116350 $D=1
M627 761 237 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=120980 $D=1
M628 550 546 760 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=116350 $D=1
M629 551 547 761 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=120980 $D=1
M630 7 550 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=116350 $D=1
M631 8 551 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=120980 $D=1
M632 762 552 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=116350 $D=1
M633 763 553 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=120980 $D=1
M634 550 548 762 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=116350 $D=1
M635 551 549 763 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=120980 $D=1
M636 7 556 554 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=116350 $D=1
M637 8 557 555 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=120980 $D=1
M638 556 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=116350 $D=1
M639 557 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=120980 $D=1
M640 764 240 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=116350 $D=1
M641 765 241 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=120980 $D=1
M642 558 554 764 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=116350 $D=1
M643 559 555 765 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=120980 $D=1
M644 7 558 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=116350 $D=1
M645 8 559 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=120980 $D=1
M646 766 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=116350 $D=1
M647 767 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=120980 $D=1
M648 558 556 766 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=116350 $D=1
M649 559 557 767 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=120980 $D=1
M650 560 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=116350 $D=1
M651 561 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=120980 $D=1
M652 562 560 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=116350 $D=1
M653 563 561 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=120980 $D=1
M654 114 113 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=116350 $D=1
M655 115 113 563 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=120980 $D=1
M656 564 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=116350 $D=1
M657 565 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=120980 $D=1
M658 566 564 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=116350 $D=1
M659 567 565 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=120980 $D=1
M660 768 116 566 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=116350 $D=1
M661 769 116 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=120980 $D=1
M662 7 111 768 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=116350 $D=1
M663 8 112 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=120980 $D=1
M664 568 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=116350 $D=1
M665 569 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=120980 $D=1
M666 570 568 566 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=116350 $D=1
M667 571 569 567 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=120980 $D=1
M668 9 117 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=116350 $D=1
M669 10 117 571 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=120980 $D=1
M670 573 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=116350 $D=1
M671 574 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=120980 $D=1
M672 7 577 575 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=116350 $D=1
M673 8 578 576 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=120980 $D=1
M674 579 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=116350 $D=1
M675 580 563 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=120980 $D=1
M676 577 579 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=116350 $D=1
M677 578 580 118 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=120980 $D=1
M678 573 562 577 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=116350 $D=1
M679 574 563 578 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=120980 $D=1
M680 581 575 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=116350 $D=1
M681 582 576 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=120980 $D=1
M682 121 581 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=116350 $D=1
M683 572 582 571 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=120980 $D=1
M684 562 575 121 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=116350 $D=1
M685 563 576 572 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=120980 $D=1
M686 583 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=116350 $D=1
M687 584 572 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=120980 $D=1
M688 585 575 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=116350 $D=1
M689 586 576 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=120980 $D=1
M690 587 585 583 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=116350 $D=1
M691 588 586 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=120980 $D=1
M692 570 575 587 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=116350 $D=1
M693 571 576 588 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=120980 $D=1
M694 589 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=116350 $D=1
M695 590 563 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=120980 $D=1
M696 7 570 589 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=116350 $D=1
M697 8 571 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=120980 $D=1
M698 591 587 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=116350 $D=1
M699 592 588 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=120980 $D=1
M700 788 562 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=116350 $D=1
M701 789 563 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=120980 $D=1
M702 593 570 788 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=116350 $D=1
M703 594 571 789 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=120980 $D=1
M704 790 562 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=116350 $D=1
M705 791 563 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=120980 $D=1
M706 595 570 790 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=116350 $D=1
M707 596 571 791 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=120980 $D=1
M708 599 562 597 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=116350 $D=1
M709 600 563 598 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=120980 $D=1
M710 597 570 599 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=116350 $D=1
M711 598 571 600 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=120980 $D=1
M712 7 595 597 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=116350 $D=1
M713 8 596 598 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=120980 $D=1
M714 601 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=116350 $D=1
M715 602 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=120980 $D=1
M716 603 601 589 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=116350 $D=1
M717 604 602 590 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=120980 $D=1
M718 593 124 603 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=116350 $D=1
M719 594 124 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=120980 $D=1
M720 605 601 591 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=116350 $D=1
M721 606 602 592 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=120980 $D=1
M722 599 124 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=116350 $D=1
M723 600 124 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=120980 $D=1
M724 607 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=116350 $D=1
M725 608 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=120980 $D=1
M726 609 607 605 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=116350 $D=1
M727 610 608 606 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=120980 $D=1
M728 603 125 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=116350 $D=1
M729 604 125 610 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=120980 $D=1
M730 11 609 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=116350 $D=1
M731 12 610 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=120980 $D=1
M732 611 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=116350 $D=1
M733 612 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=120980 $D=1
M734 613 611 127 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=116350 $D=1
M735 614 612 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=120980 $D=1
M736 129 126 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=116350 $D=1
M737 130 126 614 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=120980 $D=1
M738 615 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=116350 $D=1
M739 616 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=120980 $D=1
M740 617 615 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=116350 $D=1
M741 618 616 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=120980 $D=1
M742 133 126 617 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=116350 $D=1
M743 134 126 618 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=120980 $D=1
M744 619 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=116350 $D=1
M745 620 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=120980 $D=1
M746 136 619 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=116350 $D=1
M747 136 620 135 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=120980 $D=1
M748 137 126 136 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=116350 $D=1
M749 138 126 136 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=120980 $D=1
M750 621 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=116350 $D=1
M751 622 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=120980 $D=1
M752 623 621 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=116350 $D=1
M753 624 622 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=120980 $D=1
M754 139 126 623 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=116350 $D=1
M755 140 126 624 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=120980 $D=1
M756 625 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=116350 $D=1
M757 626 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=120980 $D=1
M758 627 625 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=116350 $D=1
M759 628 626 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=120980 $D=1
M760 141 126 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=116350 $D=1
M761 142 126 628 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=120980 $D=1
M762 7 562 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=116350 $D=1
M763 8 563 771 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=120980 $D=1
M764 130 770 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=116350 $D=1
M765 127 771 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=120980 $D=1
M766 629 143 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=116350 $D=1
M767 630 143 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=120980 $D=1
M768 144 629 130 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=116350 $D=1
M769 145 630 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=120980 $D=1
M770 613 143 144 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=116350 $D=1
M771 614 143 145 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=120980 $D=1
M772 631 146 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=116350 $D=1
M773 632 146 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=120980 $D=1
M774 147 631 144 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=116350 $D=1
M775 148 632 145 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=120980 $D=1
M776 617 146 147 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=116350 $D=1
M777 618 146 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=120980 $D=1
M778 633 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=116350 $D=1
M779 634 149 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=120980 $D=1
M780 119 633 147 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=116350 $D=1
M781 120 634 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=120980 $D=1
M782 136 149 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=116350 $D=1
M783 136 149 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=120980 $D=1
M784 635 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=116350 $D=1
M785 636 150 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=120980 $D=1
M786 151 635 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=116350 $D=1
M787 152 636 120 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=120980 $D=1
M788 623 150 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=116350 $D=1
M789 624 150 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=120980 $D=1
M790 637 153 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=116350 $D=1
M791 638 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=120980 $D=1
M792 212 637 151 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=116350 $D=1
M793 213 638 152 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=120980 $D=1
M794 627 153 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=116350 $D=1
M795 628 153 213 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=120980 $D=1
M796 639 154 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=116350 $D=1
M797 640 154 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=120980 $D=1
M798 641 639 111 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=116350 $D=1
M799 642 640 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=120980 $D=1
M800 9 154 641 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=116350 $D=1
M801 10 154 642 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=120980 $D=1
M802 792 552 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=116350 $D=1
M803 793 553 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=120980 $D=1
M804 643 641 792 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=116350 $D=1
M805 644 642 793 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=120980 $D=1
M806 647 552 645 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=116350 $D=1
M807 648 553 646 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=120980 $D=1
M808 645 641 647 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=116350 $D=1
M809 646 642 648 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=120980 $D=1
M810 7 643 645 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=116350 $D=1
M811 8 644 646 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=120980 $D=1
M812 794 155 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=116350 $D=1
M813 795 649 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=120980 $D=1
M814 772 647 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=116350 $D=1
M815 773 648 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=120980 $D=1
M816 649 772 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=116350 $D=1
M817 156 773 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=120980 $D=1
M818 650 552 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=116350 $D=1
M819 651 553 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=120980 $D=1
M820 7 652 650 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=116350 $D=1
M821 8 653 651 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=120980 $D=1
M822 652 641 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=116350 $D=1
M823 653 642 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=120980 $D=1
M824 796 650 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=116350 $D=1
M825 797 651 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=120980 $D=1
M826 654 155 796 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=116350 $D=1
M827 655 649 797 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=120980 $D=1
M828 657 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=116350 $D=1
M829 658 656 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=120980 $D=1
M830 798 654 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=116350 $D=1
M831 799 655 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=120980 $D=1
M832 656 657 798 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=116350 $D=1
M833 158 658 799 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=120980 $D=1
M834 660 659 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=116350 $D=1
M835 661 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=120980 $D=1
M836 7 664 662 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=116350 $D=1
M837 8 665 663 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=120980 $D=1
M838 666 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=116350 $D=1
M839 667 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=120980 $D=1
M840 664 666 659 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=116350 $D=1
M841 665 667 159 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=120980 $D=1
M842 660 114 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=116350 $D=1
M843 661 115 665 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=120980 $D=1
M844 668 662 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=116350 $D=1
M845 669 663 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=120980 $D=1
M846 160 668 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=116350 $D=1
M847 659 669 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=120980 $D=1
M848 114 662 160 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=116350 $D=1
M849 115 663 659 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=120980 $D=1
M850 670 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=116350 $D=1
M851 671 659 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=120980 $D=1
M852 672 662 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=116350 $D=1
M853 673 663 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=120980 $D=1
M854 214 672 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=116350 $D=1
M855 215 673 671 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=120980 $D=1
M856 7 662 214 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=116350 $D=1
M857 8 663 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=120980 $D=1
M858 674 161 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=116350 $D=1
M859 675 161 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=120980 $D=1
M860 676 674 214 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=116350 $D=1
M861 677 675 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=120980 $D=1
M862 11 161 676 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=116350 $D=1
M863 12 161 677 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=120980 $D=1
M864 678 162 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=116350 $D=1
M865 679 162 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=120980 $D=1
M866 162 678 676 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=116350 $D=1
M867 162 679 677 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=120980 $D=1
M868 7 162 162 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=116350 $D=1
M869 8 162 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=120980 $D=1
M870 680 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=116350 $D=1
M871 681 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=120980 $D=1
M872 7 680 682 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=116350 $D=1
M873 8 681 683 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=120980 $D=1
M874 684 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=116350 $D=1
M875 685 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=120980 $D=1
M876 686 680 162 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=116350 $D=1
M877 687 681 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=120980 $D=1
M878 7 686 774 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=116350 $D=1
M879 8 687 775 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=120980 $D=1
M880 688 774 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=116350 $D=1
M881 689 775 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=120980 $D=1
M882 686 682 688 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=116350 $D=1
M883 687 683 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=120980 $D=1
M884 690 110 688 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=116350 $D=1
M885 691 110 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=120980 $D=1
M886 7 694 692 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=116350 $D=1
M887 8 695 693 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=120980 $D=1
M888 694 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=116350 $D=1
M889 695 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=120980 $D=1
M890 776 690 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=116350 $D=1
M891 777 691 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=120980 $D=1
M892 696 692 776 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=116350 $D=1
M893 697 693 777 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=120980 $D=1
M894 7 696 114 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=116350 $D=1
M895 8 697 115 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=120980 $D=1
M896 778 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=116350 $D=1
M897 779 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=120980 $D=1
M898 696 694 778 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=116350 $D=1
M899 697 695 779 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=120980 $D=1
M900 188 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=117600 $D=0
M901 189 1 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=122230 $D=0
M902 190 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=117600 $D=0
M903 191 1 3 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=122230 $D=0
M904 7 188 190 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=117600 $D=0
M905 8 189 191 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=122230 $D=0
M906 192 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=117600 $D=0
M907 193 1 3 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=122230 $D=0
M908 2 188 192 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=117600 $D=0
M909 3 189 193 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=122230 $D=0
M910 194 1 2 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=117600 $D=0
M911 195 1 3 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=122230 $D=0
M912 2 188 194 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=117600 $D=0
M913 3 189 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=122230 $D=0
M914 198 4 194 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=117600 $D=0
M915 199 4 195 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=122230 $D=0
M916 196 4 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=117600 $D=0
M917 197 4 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=122230 $D=0
M918 200 4 192 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=117600 $D=0
M919 201 4 193 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=122230 $D=0
M920 190 196 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=117600 $D=0
M921 191 197 201 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=122230 $D=0
M922 202 5 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=117600 $D=0
M923 203 5 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=122230 $D=0
M924 204 5 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=117600 $D=0
M925 205 5 201 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=122230 $D=0
M926 198 202 204 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=117600 $D=0
M927 199 203 205 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=122230 $D=0
M928 206 6 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=117600 $D=0
M929 207 6 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=122230 $D=0
M930 208 6 7 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=117600 $D=0
M931 209 6 8 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=122230 $D=0
M932 9 206 208 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=117600 $D=0
M933 10 207 209 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=122230 $D=0
M934 210 6 11 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=117600 $D=0
M935 211 6 12 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=122230 $D=0
M936 212 206 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=117600 $D=0
M937 213 207 211 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=122230 $D=0
M938 216 6 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=117600 $D=0
M939 217 6 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=122230 $D=0
M940 204 206 216 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=117600 $D=0
M941 205 207 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=122230 $D=0
M942 220 13 216 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=117600 $D=0
M943 221 13 217 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=122230 $D=0
M944 218 13 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=117600 $D=0
M945 219 13 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=122230 $D=0
M946 222 13 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=117600 $D=0
M947 223 13 211 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=122230 $D=0
M948 208 218 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=117600 $D=0
M949 209 219 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=122230 $D=0
M950 224 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=117600 $D=0
M951 225 14 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=122230 $D=0
M952 226 14 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=117600 $D=0
M953 227 14 223 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=122230 $D=0
M954 220 224 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=117600 $D=0
M955 221 225 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=122230 $D=0
M956 163 15 228 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=117600 $D=0
M957 164 15 229 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=122230 $D=0
M958 230 16 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=117600 $D=0
M959 231 16 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=122230 $D=0
M960 232 228 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=117600 $D=0
M961 233 229 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=122230 $D=0
M962 163 232 698 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=117600 $D=0
M963 164 233 699 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=122230 $D=0
M964 234 698 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=117600 $D=0
M965 235 699 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=122230 $D=0
M966 232 15 234 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=117600 $D=0
M967 233 15 235 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=122230 $D=0
M968 234 230 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=117600 $D=0
M969 235 231 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=122230 $D=0
M970 240 238 234 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=117600 $D=0
M971 241 239 235 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=122230 $D=0
M972 238 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=117600 $D=0
M973 239 17 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=122230 $D=0
M974 163 18 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=117600 $D=0
M975 164 18 243 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=122230 $D=0
M976 244 19 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=117600 $D=0
M977 245 19 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=122230 $D=0
M978 246 242 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=117600 $D=0
M979 247 243 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=122230 $D=0
M980 163 246 700 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=117600 $D=0
M981 164 247 701 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=122230 $D=0
M982 248 700 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=117600 $D=0
M983 249 701 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=122230 $D=0
M984 246 18 248 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=117600 $D=0
M985 247 18 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=122230 $D=0
M986 248 244 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=117600 $D=0
M987 249 245 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=122230 $D=0
M988 240 250 248 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=117600 $D=0
M989 241 251 249 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=122230 $D=0
M990 250 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=117600 $D=0
M991 251 20 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=122230 $D=0
M992 163 21 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=117600 $D=0
M993 164 21 253 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=122230 $D=0
M994 254 22 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=117600 $D=0
M995 255 22 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=122230 $D=0
M996 256 252 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=117600 $D=0
M997 257 253 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=122230 $D=0
M998 163 256 702 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=117600 $D=0
M999 164 257 703 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=122230 $D=0
M1000 258 702 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=117600 $D=0
M1001 259 703 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=122230 $D=0
M1002 256 21 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=117600 $D=0
M1003 257 21 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=122230 $D=0
M1004 258 254 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=117600 $D=0
M1005 259 255 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=122230 $D=0
M1006 240 260 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=117600 $D=0
M1007 241 261 259 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=122230 $D=0
M1008 260 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=117600 $D=0
M1009 261 23 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=122230 $D=0
M1010 163 24 262 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=117600 $D=0
M1011 164 24 263 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=122230 $D=0
M1012 264 25 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=117600 $D=0
M1013 265 25 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=122230 $D=0
M1014 266 262 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=117600 $D=0
M1015 267 263 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=122230 $D=0
M1016 163 266 704 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=117600 $D=0
M1017 164 267 705 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=122230 $D=0
M1018 268 704 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=117600 $D=0
M1019 269 705 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=122230 $D=0
M1020 266 24 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=117600 $D=0
M1021 267 24 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=122230 $D=0
M1022 268 264 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=117600 $D=0
M1023 269 265 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=122230 $D=0
M1024 240 270 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=117600 $D=0
M1025 241 271 269 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=122230 $D=0
M1026 270 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=117600 $D=0
M1027 271 26 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=122230 $D=0
M1028 163 27 272 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=117600 $D=0
M1029 164 27 273 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=122230 $D=0
M1030 274 28 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=117600 $D=0
M1031 275 28 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=122230 $D=0
M1032 276 272 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=117600 $D=0
M1033 277 273 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=122230 $D=0
M1034 163 276 706 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=117600 $D=0
M1035 164 277 707 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=122230 $D=0
M1036 278 706 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=117600 $D=0
M1037 279 707 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=122230 $D=0
M1038 276 27 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=117600 $D=0
M1039 277 27 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=122230 $D=0
M1040 278 274 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=117600 $D=0
M1041 279 275 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=122230 $D=0
M1042 240 280 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=117600 $D=0
M1043 241 281 279 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=122230 $D=0
M1044 280 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=117600 $D=0
M1045 281 29 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=122230 $D=0
M1046 163 30 282 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=117600 $D=0
M1047 164 30 283 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=122230 $D=0
M1048 284 31 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=117600 $D=0
M1049 285 31 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=122230 $D=0
M1050 286 282 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=117600 $D=0
M1051 287 283 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=122230 $D=0
M1052 163 286 708 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=117600 $D=0
M1053 164 287 709 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=122230 $D=0
M1054 288 708 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=117600 $D=0
M1055 289 709 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=122230 $D=0
M1056 286 30 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=117600 $D=0
M1057 287 30 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=122230 $D=0
M1058 288 284 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=117600 $D=0
M1059 289 285 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=122230 $D=0
M1060 240 290 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=117600 $D=0
M1061 241 291 289 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=122230 $D=0
M1062 290 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=117600 $D=0
M1063 291 32 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=122230 $D=0
M1064 163 33 292 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=117600 $D=0
M1065 164 33 293 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=122230 $D=0
M1066 294 34 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=117600 $D=0
M1067 295 34 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=122230 $D=0
M1068 296 292 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=117600 $D=0
M1069 297 293 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=122230 $D=0
M1070 163 296 710 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=117600 $D=0
M1071 164 297 711 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=122230 $D=0
M1072 298 710 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=117600 $D=0
M1073 299 711 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=122230 $D=0
M1074 296 33 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=117600 $D=0
M1075 297 33 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=122230 $D=0
M1076 298 294 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=117600 $D=0
M1077 299 295 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=122230 $D=0
M1078 240 300 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=117600 $D=0
M1079 241 301 299 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=122230 $D=0
M1080 300 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=117600 $D=0
M1081 301 35 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=122230 $D=0
M1082 163 36 302 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=117600 $D=0
M1083 164 36 303 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=122230 $D=0
M1084 304 37 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=117600 $D=0
M1085 305 37 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=122230 $D=0
M1086 306 302 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=117600 $D=0
M1087 307 303 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=122230 $D=0
M1088 163 306 712 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=117600 $D=0
M1089 164 307 713 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=122230 $D=0
M1090 308 712 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=117600 $D=0
M1091 309 713 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=122230 $D=0
M1092 306 36 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=117600 $D=0
M1093 307 36 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=122230 $D=0
M1094 308 304 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=117600 $D=0
M1095 309 305 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=122230 $D=0
M1096 240 310 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=117600 $D=0
M1097 241 311 309 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=122230 $D=0
M1098 310 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=117600 $D=0
M1099 311 38 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=122230 $D=0
M1100 163 39 312 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=117600 $D=0
M1101 164 39 313 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=122230 $D=0
M1102 314 40 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=117600 $D=0
M1103 315 40 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=122230 $D=0
M1104 316 312 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=117600 $D=0
M1105 317 313 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=122230 $D=0
M1106 163 316 714 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=117600 $D=0
M1107 164 317 715 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=122230 $D=0
M1108 318 714 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=117600 $D=0
M1109 319 715 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=122230 $D=0
M1110 316 39 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=117600 $D=0
M1111 317 39 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=122230 $D=0
M1112 318 314 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=117600 $D=0
M1113 319 315 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=122230 $D=0
M1114 240 320 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=117600 $D=0
M1115 241 321 319 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=122230 $D=0
M1116 320 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=117600 $D=0
M1117 321 41 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=122230 $D=0
M1118 163 42 322 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=117600 $D=0
M1119 164 42 323 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=122230 $D=0
M1120 324 43 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=117600 $D=0
M1121 325 43 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=122230 $D=0
M1122 326 322 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=117600 $D=0
M1123 327 323 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=122230 $D=0
M1124 163 326 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=117600 $D=0
M1125 164 327 717 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=122230 $D=0
M1126 328 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=117600 $D=0
M1127 329 717 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=122230 $D=0
M1128 326 42 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=117600 $D=0
M1129 327 42 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=122230 $D=0
M1130 328 324 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=117600 $D=0
M1131 329 325 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=122230 $D=0
M1132 240 330 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=117600 $D=0
M1133 241 331 329 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=122230 $D=0
M1134 330 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=117600 $D=0
M1135 331 44 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=122230 $D=0
M1136 163 45 332 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=117600 $D=0
M1137 164 45 333 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=122230 $D=0
M1138 334 46 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=117600 $D=0
M1139 335 46 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=122230 $D=0
M1140 336 332 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=117600 $D=0
M1141 337 333 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=122230 $D=0
M1142 163 336 718 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=117600 $D=0
M1143 164 337 719 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=122230 $D=0
M1144 338 718 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=117600 $D=0
M1145 339 719 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=122230 $D=0
M1146 336 45 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=117600 $D=0
M1147 337 45 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=122230 $D=0
M1148 338 334 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=117600 $D=0
M1149 339 335 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=122230 $D=0
M1150 240 340 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=117600 $D=0
M1151 241 341 339 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=122230 $D=0
M1152 340 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=117600 $D=0
M1153 341 47 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=122230 $D=0
M1154 163 48 342 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=117600 $D=0
M1155 164 48 343 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=122230 $D=0
M1156 344 49 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=117600 $D=0
M1157 345 49 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=122230 $D=0
M1158 346 342 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=117600 $D=0
M1159 347 343 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=122230 $D=0
M1160 163 346 720 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=117600 $D=0
M1161 164 347 721 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=122230 $D=0
M1162 348 720 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=117600 $D=0
M1163 349 721 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=122230 $D=0
M1164 346 48 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=117600 $D=0
M1165 347 48 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=122230 $D=0
M1166 348 344 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=117600 $D=0
M1167 349 345 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=122230 $D=0
M1168 240 350 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=117600 $D=0
M1169 241 351 349 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=122230 $D=0
M1170 350 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=117600 $D=0
M1171 351 50 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=122230 $D=0
M1172 163 51 352 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=117600 $D=0
M1173 164 51 353 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=122230 $D=0
M1174 354 52 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=117600 $D=0
M1175 355 52 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=122230 $D=0
M1176 356 352 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=117600 $D=0
M1177 357 353 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=122230 $D=0
M1178 163 356 722 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=117600 $D=0
M1179 164 357 723 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=122230 $D=0
M1180 358 722 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=117600 $D=0
M1181 359 723 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=122230 $D=0
M1182 356 51 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=117600 $D=0
M1183 357 51 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=122230 $D=0
M1184 358 354 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=117600 $D=0
M1185 359 355 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=122230 $D=0
M1186 240 360 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=117600 $D=0
M1187 241 361 359 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=122230 $D=0
M1188 360 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=117600 $D=0
M1189 361 53 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=122230 $D=0
M1190 163 54 362 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=117600 $D=0
M1191 164 54 363 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=122230 $D=0
M1192 364 55 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=117600 $D=0
M1193 365 55 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=122230 $D=0
M1194 366 362 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=117600 $D=0
M1195 367 363 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=122230 $D=0
M1196 163 366 724 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=117600 $D=0
M1197 164 367 725 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=122230 $D=0
M1198 368 724 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=117600 $D=0
M1199 369 725 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=122230 $D=0
M1200 366 54 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=117600 $D=0
M1201 367 54 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=122230 $D=0
M1202 368 364 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=117600 $D=0
M1203 369 365 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=122230 $D=0
M1204 240 370 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=117600 $D=0
M1205 241 371 369 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=122230 $D=0
M1206 370 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=117600 $D=0
M1207 371 56 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=122230 $D=0
M1208 163 57 372 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=117600 $D=0
M1209 164 57 373 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=122230 $D=0
M1210 374 58 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=117600 $D=0
M1211 375 58 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=122230 $D=0
M1212 376 372 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=117600 $D=0
M1213 377 373 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=122230 $D=0
M1214 163 376 726 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=117600 $D=0
M1215 164 377 727 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=122230 $D=0
M1216 378 726 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=117600 $D=0
M1217 379 727 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=122230 $D=0
M1218 376 57 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=117600 $D=0
M1219 377 57 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=122230 $D=0
M1220 378 374 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=117600 $D=0
M1221 379 375 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=122230 $D=0
M1222 240 380 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=117600 $D=0
M1223 241 381 379 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=122230 $D=0
M1224 380 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=117600 $D=0
M1225 381 59 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=122230 $D=0
M1226 163 60 382 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=117600 $D=0
M1227 164 60 383 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=122230 $D=0
M1228 384 61 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=117600 $D=0
M1229 385 61 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=122230 $D=0
M1230 386 382 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=117600 $D=0
M1231 387 383 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=122230 $D=0
M1232 163 386 728 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=117600 $D=0
M1233 164 387 729 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=122230 $D=0
M1234 388 728 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=117600 $D=0
M1235 389 729 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=122230 $D=0
M1236 386 60 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=117600 $D=0
M1237 387 60 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=122230 $D=0
M1238 388 384 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=117600 $D=0
M1239 389 385 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=122230 $D=0
M1240 240 390 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=117600 $D=0
M1241 241 391 389 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=122230 $D=0
M1242 390 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=117600 $D=0
M1243 391 62 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=122230 $D=0
M1244 163 63 392 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=117600 $D=0
M1245 164 63 393 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=122230 $D=0
M1246 394 64 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=117600 $D=0
M1247 395 64 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=122230 $D=0
M1248 396 392 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=117600 $D=0
M1249 397 393 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=122230 $D=0
M1250 163 396 730 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=117600 $D=0
M1251 164 397 731 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=122230 $D=0
M1252 398 730 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=117600 $D=0
M1253 399 731 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=122230 $D=0
M1254 396 63 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=117600 $D=0
M1255 397 63 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=122230 $D=0
M1256 398 394 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=117600 $D=0
M1257 399 395 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=122230 $D=0
M1258 240 400 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=117600 $D=0
M1259 241 401 399 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=122230 $D=0
M1260 400 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=117600 $D=0
M1261 401 65 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=122230 $D=0
M1262 163 66 402 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=117600 $D=0
M1263 164 66 403 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=122230 $D=0
M1264 404 67 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=117600 $D=0
M1265 405 67 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=122230 $D=0
M1266 406 402 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=117600 $D=0
M1267 407 403 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=122230 $D=0
M1268 163 406 732 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=117600 $D=0
M1269 164 407 733 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=122230 $D=0
M1270 408 732 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=117600 $D=0
M1271 409 733 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=122230 $D=0
M1272 406 66 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=117600 $D=0
M1273 407 66 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=122230 $D=0
M1274 408 404 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=117600 $D=0
M1275 409 405 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=122230 $D=0
M1276 240 410 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=117600 $D=0
M1277 241 411 409 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=122230 $D=0
M1278 410 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=117600 $D=0
M1279 411 68 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=122230 $D=0
M1280 163 69 412 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=117600 $D=0
M1281 164 69 413 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=122230 $D=0
M1282 414 70 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=117600 $D=0
M1283 415 70 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=122230 $D=0
M1284 416 412 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=117600 $D=0
M1285 417 413 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=122230 $D=0
M1286 163 416 734 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=117600 $D=0
M1287 164 417 735 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=122230 $D=0
M1288 418 734 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=117600 $D=0
M1289 419 735 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=122230 $D=0
M1290 416 69 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=117600 $D=0
M1291 417 69 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=122230 $D=0
M1292 418 414 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=117600 $D=0
M1293 419 415 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=122230 $D=0
M1294 240 420 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=117600 $D=0
M1295 241 421 419 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=122230 $D=0
M1296 420 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=117600 $D=0
M1297 421 71 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=122230 $D=0
M1298 163 72 422 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=117600 $D=0
M1299 164 72 423 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=122230 $D=0
M1300 424 73 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=117600 $D=0
M1301 425 73 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=122230 $D=0
M1302 426 422 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=117600 $D=0
M1303 427 423 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=122230 $D=0
M1304 163 426 736 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=117600 $D=0
M1305 164 427 737 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=122230 $D=0
M1306 428 736 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=117600 $D=0
M1307 429 737 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=122230 $D=0
M1308 426 72 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=117600 $D=0
M1309 427 72 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=122230 $D=0
M1310 428 424 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=117600 $D=0
M1311 429 425 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=122230 $D=0
M1312 240 430 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=117600 $D=0
M1313 241 431 429 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=122230 $D=0
M1314 430 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=117600 $D=0
M1315 431 74 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=122230 $D=0
M1316 163 75 432 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=117600 $D=0
M1317 164 75 433 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=122230 $D=0
M1318 434 76 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=117600 $D=0
M1319 435 76 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=122230 $D=0
M1320 436 432 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=117600 $D=0
M1321 437 433 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=122230 $D=0
M1322 163 436 738 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=117600 $D=0
M1323 164 437 739 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=122230 $D=0
M1324 438 738 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=117600 $D=0
M1325 439 739 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=122230 $D=0
M1326 436 75 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=117600 $D=0
M1327 437 75 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=122230 $D=0
M1328 438 434 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=117600 $D=0
M1329 439 435 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=122230 $D=0
M1330 240 440 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=117600 $D=0
M1331 241 441 439 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=122230 $D=0
M1332 440 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=117600 $D=0
M1333 441 77 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=122230 $D=0
M1334 163 78 442 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=117600 $D=0
M1335 164 78 443 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=122230 $D=0
M1336 444 79 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=117600 $D=0
M1337 445 79 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=122230 $D=0
M1338 446 442 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=117600 $D=0
M1339 447 443 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=122230 $D=0
M1340 163 446 740 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=117600 $D=0
M1341 164 447 741 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=122230 $D=0
M1342 448 740 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=117600 $D=0
M1343 449 741 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=122230 $D=0
M1344 446 78 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=117600 $D=0
M1345 447 78 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=122230 $D=0
M1346 448 444 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=117600 $D=0
M1347 449 445 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=122230 $D=0
M1348 240 450 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=117600 $D=0
M1349 241 451 449 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=122230 $D=0
M1350 450 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=117600 $D=0
M1351 451 80 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=122230 $D=0
M1352 163 81 452 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=117600 $D=0
M1353 164 81 453 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=122230 $D=0
M1354 454 82 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=117600 $D=0
M1355 455 82 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=122230 $D=0
M1356 456 452 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=117600 $D=0
M1357 457 453 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=122230 $D=0
M1358 163 456 742 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=117600 $D=0
M1359 164 457 743 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=122230 $D=0
M1360 458 742 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=117600 $D=0
M1361 459 743 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=122230 $D=0
M1362 456 81 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=117600 $D=0
M1363 457 81 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=122230 $D=0
M1364 458 454 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=117600 $D=0
M1365 459 455 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=122230 $D=0
M1366 240 460 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=117600 $D=0
M1367 241 461 459 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=122230 $D=0
M1368 460 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=117600 $D=0
M1369 461 83 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=122230 $D=0
M1370 163 84 462 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=117600 $D=0
M1371 164 84 463 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=122230 $D=0
M1372 464 85 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=117600 $D=0
M1373 465 85 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=122230 $D=0
M1374 466 462 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=117600 $D=0
M1375 467 463 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=122230 $D=0
M1376 163 466 744 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=117600 $D=0
M1377 164 467 745 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=122230 $D=0
M1378 468 744 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=117600 $D=0
M1379 469 745 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=122230 $D=0
M1380 466 84 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=117600 $D=0
M1381 467 84 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=122230 $D=0
M1382 468 464 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=117600 $D=0
M1383 469 465 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=122230 $D=0
M1384 240 470 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=117600 $D=0
M1385 241 471 469 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=122230 $D=0
M1386 470 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=117600 $D=0
M1387 471 86 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=122230 $D=0
M1388 163 87 472 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=117600 $D=0
M1389 164 87 473 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=122230 $D=0
M1390 474 88 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=117600 $D=0
M1391 475 88 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=122230 $D=0
M1392 476 472 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=117600 $D=0
M1393 477 473 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=122230 $D=0
M1394 163 476 746 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=117600 $D=0
M1395 164 477 747 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=122230 $D=0
M1396 478 746 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=117600 $D=0
M1397 479 747 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=122230 $D=0
M1398 476 87 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=117600 $D=0
M1399 477 87 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=122230 $D=0
M1400 478 474 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=117600 $D=0
M1401 479 475 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=122230 $D=0
M1402 240 480 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=117600 $D=0
M1403 241 481 479 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=122230 $D=0
M1404 480 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=117600 $D=0
M1405 481 89 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=122230 $D=0
M1406 163 90 482 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=117600 $D=0
M1407 164 90 483 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=122230 $D=0
M1408 484 91 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=117600 $D=0
M1409 485 91 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=122230 $D=0
M1410 486 482 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=117600 $D=0
M1411 487 483 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=122230 $D=0
M1412 163 486 748 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=117600 $D=0
M1413 164 487 749 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=122230 $D=0
M1414 488 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=117600 $D=0
M1415 489 749 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=122230 $D=0
M1416 486 90 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=117600 $D=0
M1417 487 90 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=122230 $D=0
M1418 488 484 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=117600 $D=0
M1419 489 485 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=122230 $D=0
M1420 240 490 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=117600 $D=0
M1421 241 491 489 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=122230 $D=0
M1422 490 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=117600 $D=0
M1423 491 92 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=122230 $D=0
M1424 163 93 492 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=117600 $D=0
M1425 164 93 493 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=122230 $D=0
M1426 494 94 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=117600 $D=0
M1427 495 94 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=122230 $D=0
M1428 496 492 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=117600 $D=0
M1429 497 493 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=122230 $D=0
M1430 163 496 750 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=117600 $D=0
M1431 164 497 751 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=122230 $D=0
M1432 498 750 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=117600 $D=0
M1433 499 751 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=122230 $D=0
M1434 496 93 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=117600 $D=0
M1435 497 93 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=122230 $D=0
M1436 498 494 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=117600 $D=0
M1437 499 495 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=122230 $D=0
M1438 240 500 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=117600 $D=0
M1439 241 501 499 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=122230 $D=0
M1440 500 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=117600 $D=0
M1441 501 95 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=122230 $D=0
M1442 163 96 502 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=117600 $D=0
M1443 164 96 503 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=122230 $D=0
M1444 504 97 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=117600 $D=0
M1445 505 97 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=122230 $D=0
M1446 506 502 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=117600 $D=0
M1447 507 503 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=122230 $D=0
M1448 163 506 752 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=117600 $D=0
M1449 164 507 753 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=122230 $D=0
M1450 508 752 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=117600 $D=0
M1451 509 753 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=122230 $D=0
M1452 506 96 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=117600 $D=0
M1453 507 96 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=122230 $D=0
M1454 508 504 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=117600 $D=0
M1455 509 505 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=122230 $D=0
M1456 240 510 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=117600 $D=0
M1457 241 511 509 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=122230 $D=0
M1458 510 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=117600 $D=0
M1459 511 98 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=122230 $D=0
M1460 163 99 512 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=117600 $D=0
M1461 164 99 513 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=122230 $D=0
M1462 514 100 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=117600 $D=0
M1463 515 100 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=122230 $D=0
M1464 516 512 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=117600 $D=0
M1465 517 513 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=122230 $D=0
M1466 163 516 754 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=117600 $D=0
M1467 164 517 755 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=122230 $D=0
M1468 518 754 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=117600 $D=0
M1469 519 755 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=122230 $D=0
M1470 516 99 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=117600 $D=0
M1471 517 99 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=122230 $D=0
M1472 518 514 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=117600 $D=0
M1473 519 515 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=122230 $D=0
M1474 240 520 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=117600 $D=0
M1475 241 521 519 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=122230 $D=0
M1476 520 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=117600 $D=0
M1477 521 101 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=122230 $D=0
M1478 163 102 522 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=117600 $D=0
M1479 164 102 523 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=122230 $D=0
M1480 524 103 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=117600 $D=0
M1481 525 103 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=122230 $D=0
M1482 526 522 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=117600 $D=0
M1483 527 523 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=122230 $D=0
M1484 163 526 756 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=117600 $D=0
M1485 164 527 757 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=122230 $D=0
M1486 528 756 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=117600 $D=0
M1487 529 757 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=122230 $D=0
M1488 526 102 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=117600 $D=0
M1489 527 102 529 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=122230 $D=0
M1490 528 524 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=117600 $D=0
M1491 529 525 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=122230 $D=0
M1492 240 530 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=117600 $D=0
M1493 241 531 529 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=122230 $D=0
M1494 530 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=117600 $D=0
M1495 531 104 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=122230 $D=0
M1496 163 105 532 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=117600 $D=0
M1497 164 105 533 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=122230 $D=0
M1498 534 106 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=117600 $D=0
M1499 535 106 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=122230 $D=0
M1500 536 532 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=117600 $D=0
M1501 537 533 227 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=122230 $D=0
M1502 163 536 758 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=117600 $D=0
M1503 164 537 759 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=122230 $D=0
M1504 538 758 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=117600 $D=0
M1505 539 759 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=122230 $D=0
M1506 536 105 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=117600 $D=0
M1507 537 105 539 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=122230 $D=0
M1508 538 534 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=117600 $D=0
M1509 539 535 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=122230 $D=0
M1510 240 540 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=117600 $D=0
M1511 241 541 539 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=122230 $D=0
M1512 540 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=117600 $D=0
M1513 541 107 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=122230 $D=0
M1514 163 108 542 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=117600 $D=0
M1515 164 108 543 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=122230 $D=0
M1516 544 109 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=117600 $D=0
M1517 545 109 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=122230 $D=0
M1518 7 544 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=117600 $D=0
M1519 8 545 237 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=122230 $D=0
M1520 240 542 7 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=117600 $D=0
M1521 241 543 8 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=122230 $D=0
M1522 163 548 546 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=117600 $D=0
M1523 164 549 547 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=122230 $D=0
M1524 548 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=117600 $D=0
M1525 549 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=122230 $D=0
M1526 760 236 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=117600 $D=0
M1527 761 237 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=122230 $D=0
M1528 550 548 760 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=117600 $D=0
M1529 551 549 761 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=122230 $D=0
M1530 163 550 552 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=117600 $D=0
M1531 164 551 553 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=122230 $D=0
M1532 762 552 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=117600 $D=0
M1533 763 553 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=122230 $D=0
M1534 550 546 762 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=117600 $D=0
M1535 551 547 763 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=122230 $D=0
M1536 163 556 554 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=117600 $D=0
M1537 164 557 555 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=122230 $D=0
M1538 556 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=117600 $D=0
M1539 557 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=122230 $D=0
M1540 764 240 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=117600 $D=0
M1541 765 241 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=122230 $D=0
M1542 558 556 764 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=117600 $D=0
M1543 559 557 765 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=122230 $D=0
M1544 163 558 111 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=117600 $D=0
M1545 164 559 112 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=122230 $D=0
M1546 766 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=117600 $D=0
M1547 767 112 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=122230 $D=0
M1548 558 554 766 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=117600 $D=0
M1549 559 555 767 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=122230 $D=0
M1550 560 113 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=117600 $D=0
M1551 561 113 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=122230 $D=0
M1552 562 113 552 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=117600 $D=0
M1553 563 113 553 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=122230 $D=0
M1554 114 560 562 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=117600 $D=0
M1555 115 561 563 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=122230 $D=0
M1556 564 116 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=117600 $D=0
M1557 565 116 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=122230 $D=0
M1558 566 116 111 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=117600 $D=0
M1559 567 116 112 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=122230 $D=0
M1560 768 564 566 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=117600 $D=0
M1561 769 565 567 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=122230 $D=0
M1562 163 111 768 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=117600 $D=0
M1563 164 112 769 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=122230 $D=0
M1564 568 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=117600 $D=0
M1565 569 117 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=122230 $D=0
M1566 570 117 566 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=117600 $D=0
M1567 571 117 567 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=122230 $D=0
M1568 9 568 570 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=117600 $D=0
M1569 10 569 571 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=122230 $D=0
M1570 573 572 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=117600 $D=0
M1571 574 118 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=122230 $D=0
M1572 163 577 575 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=117600 $D=0
M1573 164 578 576 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=122230 $D=0
M1574 579 562 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=117600 $D=0
M1575 580 563 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=122230 $D=0
M1576 577 562 572 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=117600 $D=0
M1577 578 563 118 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=122230 $D=0
M1578 573 579 577 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=117600 $D=0
M1579 574 580 578 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=122230 $D=0
M1580 581 575 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=117600 $D=0
M1581 582 576 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=122230 $D=0
M1582 121 575 570 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=117600 $D=0
M1583 572 576 571 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=122230 $D=0
M1584 562 581 121 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=117600 $D=0
M1585 563 582 572 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=122230 $D=0
M1586 583 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=117600 $D=0
M1587 584 572 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=122230 $D=0
M1588 585 575 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=117600 $D=0
M1589 586 576 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=122230 $D=0
M1590 587 575 583 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=117600 $D=0
M1591 588 576 584 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=122230 $D=0
M1592 570 585 587 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=117600 $D=0
M1593 571 586 588 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=122230 $D=0
M1594 780 562 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=117240 $D=0
M1595 781 563 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=121870 $D=0
M1596 589 570 780 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=117240 $D=0
M1597 590 571 781 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=121870 $D=0
M1598 591 587 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=117600 $D=0
M1599 592 588 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=122230 $D=0
M1600 593 562 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=117600 $D=0
M1601 594 563 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=122230 $D=0
M1602 163 570 593 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=117600 $D=0
M1603 164 571 594 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=122230 $D=0
M1604 595 562 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=117600 $D=0
M1605 596 563 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=122230 $D=0
M1606 163 570 595 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=117600 $D=0
M1607 164 571 596 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=122230 $D=0
M1608 782 562 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=117420 $D=0
M1609 783 563 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=122050 $D=0
M1610 599 570 782 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=117420 $D=0
M1611 600 571 783 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=122050 $D=0
M1612 163 595 599 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=117600 $D=0
M1613 164 596 600 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=122230 $D=0
M1614 601 124 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=117600 $D=0
M1615 602 124 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=122230 $D=0
M1616 603 124 589 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=117600 $D=0
M1617 604 124 590 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=122230 $D=0
M1618 593 601 603 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=117600 $D=0
M1619 594 602 604 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=122230 $D=0
M1620 605 124 591 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=117600 $D=0
M1621 606 124 592 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=122230 $D=0
M1622 599 601 605 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=117600 $D=0
M1623 600 602 606 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=122230 $D=0
M1624 607 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=117600 $D=0
M1625 608 125 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=122230 $D=0
M1626 609 125 605 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=117600 $D=0
M1627 610 125 606 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=122230 $D=0
M1628 603 607 609 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=117600 $D=0
M1629 604 608 610 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=122230 $D=0
M1630 11 609 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=117600 $D=0
M1631 12 610 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=122230 $D=0
M1632 611 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=117600 $D=0
M1633 612 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=122230 $D=0
M1634 613 126 127 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=117600 $D=0
M1635 614 126 128 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=122230 $D=0
M1636 129 611 613 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=117600 $D=0
M1637 130 612 614 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=122230 $D=0
M1638 615 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=117600 $D=0
M1639 616 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=122230 $D=0
M1640 617 126 131 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=117600 $D=0
M1641 618 126 132 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=122230 $D=0
M1642 133 615 617 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=117600 $D=0
M1643 134 616 618 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=122230 $D=0
M1644 619 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=117600 $D=0
M1645 620 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=122230 $D=0
M1646 136 126 122 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=117600 $D=0
M1647 136 126 135 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=122230 $D=0
M1648 137 619 136 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=117600 $D=0
M1649 138 620 136 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=122230 $D=0
M1650 621 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=117600 $D=0
M1651 622 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=122230 $D=0
M1652 623 126 7 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=117600 $D=0
M1653 624 126 8 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=122230 $D=0
M1654 139 621 623 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=117600 $D=0
M1655 140 622 624 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=122230 $D=0
M1656 625 126 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=117600 $D=0
M1657 626 126 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=122230 $D=0
M1658 627 126 7 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=117600 $D=0
M1659 628 126 8 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=122230 $D=0
M1660 141 625 627 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=117600 $D=0
M1661 142 626 628 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=122230 $D=0
M1662 163 562 770 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=117600 $D=0
M1663 164 563 771 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=122230 $D=0
M1664 130 770 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=117600 $D=0
M1665 127 771 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=122230 $D=0
M1666 629 143 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=117600 $D=0
M1667 630 143 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=122230 $D=0
M1668 144 143 130 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=117600 $D=0
M1669 145 143 127 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=122230 $D=0
M1670 613 629 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=117600 $D=0
M1671 614 630 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=122230 $D=0
M1672 631 146 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=117600 $D=0
M1673 632 146 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=122230 $D=0
M1674 147 146 144 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=117600 $D=0
M1675 148 146 145 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=122230 $D=0
M1676 617 631 147 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=117600 $D=0
M1677 618 632 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=122230 $D=0
M1678 633 149 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=117600 $D=0
M1679 634 149 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=122230 $D=0
M1680 119 149 147 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=117600 $D=0
M1681 120 149 148 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=122230 $D=0
M1682 136 633 119 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=117600 $D=0
M1683 136 634 120 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=122230 $D=0
M1684 635 150 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=117600 $D=0
M1685 636 150 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=122230 $D=0
M1686 151 150 119 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=117600 $D=0
M1687 152 150 120 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=122230 $D=0
M1688 623 635 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=117600 $D=0
M1689 624 636 152 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=122230 $D=0
M1690 637 153 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=117600 $D=0
M1691 638 153 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=122230 $D=0
M1692 212 153 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=117600 $D=0
M1693 213 153 152 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=122230 $D=0
M1694 627 637 212 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=117600 $D=0
M1695 628 638 213 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=122230 $D=0
M1696 639 154 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=117600 $D=0
M1697 640 154 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=122230 $D=0
M1698 641 154 111 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=117600 $D=0
M1699 642 154 112 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=122230 $D=0
M1700 9 639 641 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=117600 $D=0
M1701 10 640 642 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=122230 $D=0
M1702 643 552 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=117600 $D=0
M1703 644 553 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=122230 $D=0
M1704 163 641 643 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=117600 $D=0
M1705 164 642 644 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=122230 $D=0
M1706 784 552 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=117420 $D=0
M1707 785 553 164 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=122050 $D=0
M1708 647 641 784 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=117420 $D=0
M1709 648 642 785 164 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=122050 $D=0
M1710 163 643 647 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=117600 $D=0
M1711 164 644 648 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=122230 $D=0
M1712 772 155 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=117600 $D=0
M1713 773 649 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=122230 $D=0
M1714 163 647 772 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=117600 $D=0
M1715 164 648 773 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=122230 $D=0
M1716 649 772 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=117600 $D=0
M1717 156 773 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=122230 $D=0
M1718 786 552 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=117240 $D=0
M1719 787 553 164 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=121870 $D=0
M1720 650 652 786 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=117240 $D=0
M1721 651 653 787 164 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=121870 $D=0
M1722 652 641 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=117600 $D=0
M1723 653 642 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=122230 $D=0
M1724 654 650 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=117600 $D=0
M1725 655 651 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=122230 $D=0
M1726 163 155 654 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=117600 $D=0
M1727 164 649 655 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=122230 $D=0
M1728 657 157 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=117600 $D=0
M1729 658 656 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=122230 $D=0
M1730 656 654 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=117600 $D=0
M1731 158 655 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=122230 $D=0
M1732 163 657 656 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=117600 $D=0
M1733 164 658 158 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=122230 $D=0
M1734 660 659 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=117600 $D=0
M1735 661 159 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=122230 $D=0
M1736 163 664 662 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=117600 $D=0
M1737 164 665 663 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=122230 $D=0
M1738 666 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=117600 $D=0
M1739 667 115 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=122230 $D=0
M1740 664 114 659 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=117600 $D=0
M1741 665 115 159 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=122230 $D=0
M1742 660 666 664 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=117600 $D=0
M1743 661 667 665 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=122230 $D=0
M1744 668 662 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=117600 $D=0
M1745 669 663 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=122230 $D=0
M1746 160 662 7 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=117600 $D=0
M1747 659 663 8 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=122230 $D=0
M1748 114 668 160 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=117600 $D=0
M1749 115 669 659 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=122230 $D=0
M1750 670 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=117600 $D=0
M1751 671 659 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=122230 $D=0
M1752 672 662 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=117600 $D=0
M1753 673 663 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=122230 $D=0
M1754 214 662 670 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=117600 $D=0
M1755 215 663 671 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=122230 $D=0
M1756 7 672 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=117600 $D=0
M1757 8 673 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=122230 $D=0
M1758 674 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=117600 $D=0
M1759 675 161 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=122230 $D=0
M1760 676 161 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=117600 $D=0
M1761 677 161 215 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=122230 $D=0
M1762 11 674 676 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=117600 $D=0
M1763 12 675 677 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=122230 $D=0
M1764 678 162 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=117600 $D=0
M1765 679 162 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=122230 $D=0
M1766 162 162 676 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=117600 $D=0
M1767 162 162 677 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=122230 $D=0
M1768 7 678 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=117600 $D=0
M1769 8 679 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=122230 $D=0
M1770 680 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=117600 $D=0
M1771 681 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=122230 $D=0
M1772 163 680 682 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=117600 $D=0
M1773 164 681 683 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=122230 $D=0
M1774 684 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=117600 $D=0
M1775 685 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=122230 $D=0
M1776 686 682 162 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=117600 $D=0
M1777 687 683 162 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=122230 $D=0
M1778 163 686 774 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=117600 $D=0
M1779 164 687 775 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=122230 $D=0
M1780 688 774 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=117600 $D=0
M1781 689 775 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=122230 $D=0
M1782 686 680 688 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=117600 $D=0
M1783 687 681 689 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=122230 $D=0
M1784 690 684 688 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=117600 $D=0
M1785 691 685 689 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=122230 $D=0
M1786 163 694 692 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=117600 $D=0
M1787 164 695 693 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=122230 $D=0
M1788 694 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=117600 $D=0
M1789 695 110 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=122230 $D=0
M1790 776 690 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=117600 $D=0
M1791 777 691 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=122230 $D=0
M1792 696 694 776 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=117600 $D=0
M1793 697 695 777 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=122230 $D=0
M1794 163 696 114 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=117600 $D=0
M1795 164 697 115 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=122230 $D=0
M1796 778 114 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=117600 $D=0
M1797 779 115 164 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=122230 $D=0
M1798 696 692 778 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=117600 $D=0
M1799 697 693 779 164 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=122230 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162
** N=806 EP=162 IP=1514 FDC=1800
M0 194 1 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=107090 $D=1
M1 195 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=111720 $D=1
M2 196 194 2 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=107090 $D=1
M3 197 195 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=111720 $D=1
M4 4 1 196 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=107090 $D=1
M5 8 1 197 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=111720 $D=1
M6 198 194 3 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=107090 $D=1
M7 199 195 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=111720 $D=1
M8 2 1 198 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=107090 $D=1
M9 3 1 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=111720 $D=1
M10 200 194 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=107090 $D=1
M11 201 195 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=111720 $D=1
M12 2 1 200 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=107090 $D=1
M13 3 1 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=111720 $D=1
M14 204 202 200 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=107090 $D=1
M15 205 203 201 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=111720 $D=1
M16 202 5 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=107090 $D=1
M17 203 5 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=111720 $D=1
M18 206 202 198 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=107090 $D=1
M19 207 203 199 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=111720 $D=1
M20 196 5 206 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=107090 $D=1
M21 197 5 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=111720 $D=1
M22 208 6 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=107090 $D=1
M23 209 6 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=111720 $D=1
M24 210 208 206 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=107090 $D=1
M25 211 209 207 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=111720 $D=1
M26 204 6 210 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=107090 $D=1
M27 205 6 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=111720 $D=1
M28 212 7 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=107090 $D=1
M29 213 7 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=111720 $D=1
M30 214 212 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=107090 $D=1
M31 215 213 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=111720 $D=1
M32 9 7 214 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=107090 $D=1
M33 10 7 215 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=111720 $D=1
M34 216 212 11 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=107090 $D=1
M35 217 213 12 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=111720 $D=1
M36 218 7 216 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=107090 $D=1
M37 219 7 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=111720 $D=1
M38 222 212 220 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=107090 $D=1
M39 223 213 221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=111720 $D=1
M40 210 7 222 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=107090 $D=1
M41 211 7 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=111720 $D=1
M42 226 224 222 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=107090 $D=1
M43 227 225 223 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=111720 $D=1
M44 224 13 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=107090 $D=1
M45 225 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=111720 $D=1
M46 228 224 216 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=107090 $D=1
M47 229 225 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=111720 $D=1
M48 214 13 228 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=107090 $D=1
M49 215 13 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=111720 $D=1
M50 230 14 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=107090 $D=1
M51 231 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=111720 $D=1
M52 232 230 228 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=107090 $D=1
M53 233 231 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=111720 $D=1
M54 226 14 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=107090 $D=1
M55 227 14 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=111720 $D=1
M56 4 15 234 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=107090 $D=1
M57 8 15 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=111720 $D=1
M58 236 16 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=107090 $D=1
M59 237 16 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=111720 $D=1
M60 238 15 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=107090 $D=1
M61 239 15 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=111720 $D=1
M62 4 238 705 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=107090 $D=1
M63 8 239 706 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=111720 $D=1
M64 240 705 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=107090 $D=1
M65 241 706 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=111720 $D=1
M66 238 234 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=107090 $D=1
M67 239 235 241 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=111720 $D=1
M68 240 16 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=107090 $D=1
M69 241 16 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=111720 $D=1
M70 246 17 240 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=107090 $D=1
M71 247 17 241 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=111720 $D=1
M72 244 17 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=107090 $D=1
M73 245 17 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=111720 $D=1
M74 4 18 248 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=107090 $D=1
M75 8 18 249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=111720 $D=1
M76 250 19 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=107090 $D=1
M77 251 19 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=111720 $D=1
M78 252 18 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=107090 $D=1
M79 253 18 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=111720 $D=1
M80 4 252 707 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=107090 $D=1
M81 8 253 708 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=111720 $D=1
M82 254 707 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=107090 $D=1
M83 255 708 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=111720 $D=1
M84 252 248 254 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=107090 $D=1
M85 253 249 255 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=111720 $D=1
M86 254 19 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=107090 $D=1
M87 255 19 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=111720 $D=1
M88 246 20 254 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=107090 $D=1
M89 247 20 255 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=111720 $D=1
M90 256 20 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=107090 $D=1
M91 257 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=111720 $D=1
M92 4 21 258 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=107090 $D=1
M93 8 21 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=111720 $D=1
M94 260 22 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=107090 $D=1
M95 261 22 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=111720 $D=1
M96 262 21 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=107090 $D=1
M97 263 21 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=111720 $D=1
M98 4 262 709 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=107090 $D=1
M99 8 263 710 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=111720 $D=1
M100 264 709 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=107090 $D=1
M101 265 710 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=111720 $D=1
M102 262 258 264 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=107090 $D=1
M103 263 259 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=111720 $D=1
M104 264 22 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=107090 $D=1
M105 265 22 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=111720 $D=1
M106 246 23 264 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=107090 $D=1
M107 247 23 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=111720 $D=1
M108 266 23 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=107090 $D=1
M109 267 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=111720 $D=1
M110 4 24 268 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=107090 $D=1
M111 8 24 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=111720 $D=1
M112 270 25 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=107090 $D=1
M113 271 25 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=111720 $D=1
M114 272 24 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=107090 $D=1
M115 273 24 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=111720 $D=1
M116 4 272 711 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=107090 $D=1
M117 8 273 712 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=111720 $D=1
M118 274 711 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=107090 $D=1
M119 275 712 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=111720 $D=1
M120 272 268 274 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=107090 $D=1
M121 273 269 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=111720 $D=1
M122 274 25 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=107090 $D=1
M123 275 25 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=111720 $D=1
M124 246 26 274 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=107090 $D=1
M125 247 26 275 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=111720 $D=1
M126 276 26 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=107090 $D=1
M127 277 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=111720 $D=1
M128 4 27 278 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=107090 $D=1
M129 8 27 279 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=111720 $D=1
M130 280 28 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=107090 $D=1
M131 281 28 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=111720 $D=1
M132 282 27 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=107090 $D=1
M133 283 27 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=111720 $D=1
M134 4 282 713 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=107090 $D=1
M135 8 283 714 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=111720 $D=1
M136 284 713 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=107090 $D=1
M137 285 714 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=111720 $D=1
M138 282 278 284 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=107090 $D=1
M139 283 279 285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=111720 $D=1
M140 284 28 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=107090 $D=1
M141 285 28 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=111720 $D=1
M142 246 29 284 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=107090 $D=1
M143 247 29 285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=111720 $D=1
M144 286 29 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=107090 $D=1
M145 287 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=111720 $D=1
M146 4 30 288 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=107090 $D=1
M147 8 30 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=111720 $D=1
M148 290 31 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=107090 $D=1
M149 291 31 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=111720 $D=1
M150 292 30 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=107090 $D=1
M151 293 30 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=111720 $D=1
M152 4 292 715 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=107090 $D=1
M153 8 293 716 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=111720 $D=1
M154 294 715 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=107090 $D=1
M155 295 716 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=111720 $D=1
M156 292 288 294 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=107090 $D=1
M157 293 289 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=111720 $D=1
M158 294 31 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=107090 $D=1
M159 295 31 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=111720 $D=1
M160 246 32 294 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=107090 $D=1
M161 247 32 295 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=111720 $D=1
M162 296 32 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=107090 $D=1
M163 297 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=111720 $D=1
M164 4 33 298 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=107090 $D=1
M165 8 33 299 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=111720 $D=1
M166 300 34 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=107090 $D=1
M167 301 34 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=111720 $D=1
M168 302 33 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=107090 $D=1
M169 303 33 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=111720 $D=1
M170 4 302 717 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=107090 $D=1
M171 8 303 718 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=111720 $D=1
M172 304 717 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=107090 $D=1
M173 305 718 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=111720 $D=1
M174 302 298 304 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=107090 $D=1
M175 303 299 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=111720 $D=1
M176 304 34 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=107090 $D=1
M177 305 34 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=111720 $D=1
M178 246 35 304 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=107090 $D=1
M179 247 35 305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=111720 $D=1
M180 306 35 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=107090 $D=1
M181 307 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=111720 $D=1
M182 4 36 308 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=107090 $D=1
M183 8 36 309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=111720 $D=1
M184 310 37 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=107090 $D=1
M185 311 37 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=111720 $D=1
M186 312 36 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=107090 $D=1
M187 313 36 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=111720 $D=1
M188 4 312 719 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=107090 $D=1
M189 8 313 720 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=111720 $D=1
M190 314 719 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=107090 $D=1
M191 315 720 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=111720 $D=1
M192 312 308 314 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=107090 $D=1
M193 313 309 315 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=111720 $D=1
M194 314 37 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=107090 $D=1
M195 315 37 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=111720 $D=1
M196 246 38 314 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=107090 $D=1
M197 247 38 315 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=111720 $D=1
M198 316 38 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=107090 $D=1
M199 317 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=111720 $D=1
M200 4 39 318 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=107090 $D=1
M201 8 39 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=111720 $D=1
M202 320 40 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=107090 $D=1
M203 321 40 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=111720 $D=1
M204 322 39 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=107090 $D=1
M205 323 39 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=111720 $D=1
M206 4 322 721 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=107090 $D=1
M207 8 323 722 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=111720 $D=1
M208 324 721 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=107090 $D=1
M209 325 722 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=111720 $D=1
M210 322 318 324 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=107090 $D=1
M211 323 319 325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=111720 $D=1
M212 324 40 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=107090 $D=1
M213 325 40 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=111720 $D=1
M214 246 41 324 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=107090 $D=1
M215 247 41 325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=111720 $D=1
M216 326 41 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=107090 $D=1
M217 327 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=111720 $D=1
M218 4 42 328 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=107090 $D=1
M219 8 42 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=111720 $D=1
M220 330 43 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=107090 $D=1
M221 331 43 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=111720 $D=1
M222 332 42 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=107090 $D=1
M223 333 42 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=111720 $D=1
M224 4 332 723 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=107090 $D=1
M225 8 333 724 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=111720 $D=1
M226 334 723 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=107090 $D=1
M227 335 724 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=111720 $D=1
M228 332 328 334 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=107090 $D=1
M229 333 329 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=111720 $D=1
M230 334 43 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=107090 $D=1
M231 335 43 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=111720 $D=1
M232 246 44 334 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=107090 $D=1
M233 247 44 335 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=111720 $D=1
M234 336 44 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=107090 $D=1
M235 337 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=111720 $D=1
M236 4 45 338 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=107090 $D=1
M237 8 45 339 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=111720 $D=1
M238 340 46 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=107090 $D=1
M239 341 46 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=111720 $D=1
M240 342 45 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=107090 $D=1
M241 343 45 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=111720 $D=1
M242 4 342 725 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=107090 $D=1
M243 8 343 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=111720 $D=1
M244 344 725 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=107090 $D=1
M245 345 726 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=111720 $D=1
M246 342 338 344 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=107090 $D=1
M247 343 339 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=111720 $D=1
M248 344 46 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=107090 $D=1
M249 345 46 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=111720 $D=1
M250 246 47 344 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=107090 $D=1
M251 247 47 345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=111720 $D=1
M252 346 47 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=107090 $D=1
M253 347 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=111720 $D=1
M254 4 48 348 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=107090 $D=1
M255 8 48 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=111720 $D=1
M256 350 49 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=107090 $D=1
M257 351 49 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=111720 $D=1
M258 352 48 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=107090 $D=1
M259 353 48 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=111720 $D=1
M260 4 352 727 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=107090 $D=1
M261 8 353 728 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=111720 $D=1
M262 354 727 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=107090 $D=1
M263 355 728 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=111720 $D=1
M264 352 348 354 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=107090 $D=1
M265 353 349 355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=111720 $D=1
M266 354 49 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=107090 $D=1
M267 355 49 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=111720 $D=1
M268 246 50 354 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=107090 $D=1
M269 247 50 355 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=111720 $D=1
M270 356 50 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=107090 $D=1
M271 357 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=111720 $D=1
M272 4 51 358 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=107090 $D=1
M273 8 51 359 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=111720 $D=1
M274 360 52 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=107090 $D=1
M275 361 52 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=111720 $D=1
M276 362 51 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=107090 $D=1
M277 363 51 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=111720 $D=1
M278 4 362 729 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=107090 $D=1
M279 8 363 730 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=111720 $D=1
M280 364 729 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=107090 $D=1
M281 365 730 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=111720 $D=1
M282 362 358 364 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=107090 $D=1
M283 363 359 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=111720 $D=1
M284 364 52 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=107090 $D=1
M285 365 52 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=111720 $D=1
M286 246 53 364 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=107090 $D=1
M287 247 53 365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=111720 $D=1
M288 366 53 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=107090 $D=1
M289 367 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=111720 $D=1
M290 4 54 368 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=107090 $D=1
M291 8 54 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=111720 $D=1
M292 370 55 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=107090 $D=1
M293 371 55 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=111720 $D=1
M294 372 54 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=107090 $D=1
M295 373 54 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=111720 $D=1
M296 4 372 731 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=107090 $D=1
M297 8 373 732 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=111720 $D=1
M298 374 731 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=107090 $D=1
M299 375 732 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=111720 $D=1
M300 372 368 374 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=107090 $D=1
M301 373 369 375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=111720 $D=1
M302 374 55 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=107090 $D=1
M303 375 55 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=111720 $D=1
M304 246 56 374 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=107090 $D=1
M305 247 56 375 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=111720 $D=1
M306 376 56 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=107090 $D=1
M307 377 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=111720 $D=1
M308 4 57 378 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=107090 $D=1
M309 8 57 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=111720 $D=1
M310 380 58 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=107090 $D=1
M311 381 58 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=111720 $D=1
M312 382 57 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=107090 $D=1
M313 383 57 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=111720 $D=1
M314 4 382 733 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=107090 $D=1
M315 8 383 734 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=111720 $D=1
M316 384 733 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=107090 $D=1
M317 385 734 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=111720 $D=1
M318 382 378 384 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=107090 $D=1
M319 383 379 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=111720 $D=1
M320 384 58 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=107090 $D=1
M321 385 58 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=111720 $D=1
M322 246 59 384 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=107090 $D=1
M323 247 59 385 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=111720 $D=1
M324 386 59 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=107090 $D=1
M325 387 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=111720 $D=1
M326 4 60 388 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=107090 $D=1
M327 8 60 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=111720 $D=1
M328 390 61 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=107090 $D=1
M329 391 61 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=111720 $D=1
M330 392 60 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=107090 $D=1
M331 393 60 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=111720 $D=1
M332 4 392 735 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=107090 $D=1
M333 8 393 736 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=111720 $D=1
M334 394 735 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=107090 $D=1
M335 395 736 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=111720 $D=1
M336 392 388 394 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=107090 $D=1
M337 393 389 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=111720 $D=1
M338 394 61 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=107090 $D=1
M339 395 61 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=111720 $D=1
M340 246 62 394 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=107090 $D=1
M341 247 62 395 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=111720 $D=1
M342 396 62 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=107090 $D=1
M343 397 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=111720 $D=1
M344 4 63 398 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=107090 $D=1
M345 8 63 399 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=111720 $D=1
M346 400 64 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=107090 $D=1
M347 401 64 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=111720 $D=1
M348 402 63 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=107090 $D=1
M349 403 63 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=111720 $D=1
M350 4 402 737 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=107090 $D=1
M351 8 403 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=111720 $D=1
M352 404 737 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=107090 $D=1
M353 405 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=111720 $D=1
M354 402 398 404 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=107090 $D=1
M355 403 399 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=111720 $D=1
M356 404 64 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=107090 $D=1
M357 405 64 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=111720 $D=1
M358 246 65 404 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=107090 $D=1
M359 247 65 405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=111720 $D=1
M360 406 65 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=107090 $D=1
M361 407 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=111720 $D=1
M362 4 66 408 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=107090 $D=1
M363 8 66 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=111720 $D=1
M364 410 67 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=107090 $D=1
M365 411 67 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=111720 $D=1
M366 412 66 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=107090 $D=1
M367 413 66 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=111720 $D=1
M368 4 412 739 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=107090 $D=1
M369 8 413 740 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=111720 $D=1
M370 414 739 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=107090 $D=1
M371 415 740 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=111720 $D=1
M372 412 408 414 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=107090 $D=1
M373 413 409 415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=111720 $D=1
M374 414 67 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=107090 $D=1
M375 415 67 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=111720 $D=1
M376 246 68 414 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=107090 $D=1
M377 247 68 415 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=111720 $D=1
M378 416 68 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=107090 $D=1
M379 417 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=111720 $D=1
M380 4 69 418 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=107090 $D=1
M381 8 69 419 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=111720 $D=1
M382 420 70 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=107090 $D=1
M383 421 70 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=111720 $D=1
M384 422 69 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=107090 $D=1
M385 423 69 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=111720 $D=1
M386 4 422 741 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=107090 $D=1
M387 8 423 742 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=111720 $D=1
M388 424 741 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=107090 $D=1
M389 425 742 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=111720 $D=1
M390 422 418 424 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=107090 $D=1
M391 423 419 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=111720 $D=1
M392 424 70 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=107090 $D=1
M393 425 70 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=111720 $D=1
M394 246 71 424 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=107090 $D=1
M395 247 71 425 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=111720 $D=1
M396 426 71 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=107090 $D=1
M397 427 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=111720 $D=1
M398 4 72 428 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=107090 $D=1
M399 8 72 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=111720 $D=1
M400 430 73 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=107090 $D=1
M401 431 73 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=111720 $D=1
M402 432 72 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=107090 $D=1
M403 433 72 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=111720 $D=1
M404 4 432 743 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=107090 $D=1
M405 8 433 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=111720 $D=1
M406 434 743 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=107090 $D=1
M407 435 744 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=111720 $D=1
M408 432 428 434 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=107090 $D=1
M409 433 429 435 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=111720 $D=1
M410 434 73 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=107090 $D=1
M411 435 73 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=111720 $D=1
M412 246 74 434 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=107090 $D=1
M413 247 74 435 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=111720 $D=1
M414 436 74 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=107090 $D=1
M415 437 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=111720 $D=1
M416 4 75 438 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=107090 $D=1
M417 8 75 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=111720 $D=1
M418 440 76 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=107090 $D=1
M419 441 76 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=111720 $D=1
M420 442 75 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=107090 $D=1
M421 443 75 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=111720 $D=1
M422 4 442 745 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=107090 $D=1
M423 8 443 746 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=111720 $D=1
M424 444 745 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=107090 $D=1
M425 445 746 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=111720 $D=1
M426 442 438 444 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=107090 $D=1
M427 443 439 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=111720 $D=1
M428 444 76 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=107090 $D=1
M429 445 76 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=111720 $D=1
M430 246 77 444 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=107090 $D=1
M431 247 77 445 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=111720 $D=1
M432 446 77 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=107090 $D=1
M433 447 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=111720 $D=1
M434 4 78 448 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=107090 $D=1
M435 8 78 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=111720 $D=1
M436 450 79 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=107090 $D=1
M437 451 79 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=111720 $D=1
M438 452 78 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=107090 $D=1
M439 453 78 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=111720 $D=1
M440 4 452 747 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=107090 $D=1
M441 8 453 748 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=111720 $D=1
M442 454 747 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=107090 $D=1
M443 455 748 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=111720 $D=1
M444 452 448 454 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=107090 $D=1
M445 453 449 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=111720 $D=1
M446 454 79 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=107090 $D=1
M447 455 79 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=111720 $D=1
M448 246 80 454 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=107090 $D=1
M449 247 80 455 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=111720 $D=1
M450 456 80 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=107090 $D=1
M451 457 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=111720 $D=1
M452 4 81 458 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=107090 $D=1
M453 8 81 459 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=111720 $D=1
M454 460 82 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=107090 $D=1
M455 461 82 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=111720 $D=1
M456 462 81 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=107090 $D=1
M457 463 81 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=111720 $D=1
M458 4 462 749 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=107090 $D=1
M459 8 463 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=111720 $D=1
M460 464 749 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=107090 $D=1
M461 465 750 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=111720 $D=1
M462 462 458 464 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=107090 $D=1
M463 463 459 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=111720 $D=1
M464 464 82 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=107090 $D=1
M465 465 82 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=111720 $D=1
M466 246 83 464 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=107090 $D=1
M467 247 83 465 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=111720 $D=1
M468 466 83 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=107090 $D=1
M469 467 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=111720 $D=1
M470 4 84 468 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=107090 $D=1
M471 8 84 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=111720 $D=1
M472 470 85 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=107090 $D=1
M473 471 85 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=111720 $D=1
M474 472 84 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=107090 $D=1
M475 473 84 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=111720 $D=1
M476 4 472 751 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=107090 $D=1
M477 8 473 752 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=111720 $D=1
M478 474 751 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=107090 $D=1
M479 475 752 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=111720 $D=1
M480 472 468 474 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=107090 $D=1
M481 473 469 475 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=111720 $D=1
M482 474 85 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=107090 $D=1
M483 475 85 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=111720 $D=1
M484 246 86 474 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=107090 $D=1
M485 247 86 475 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=111720 $D=1
M486 476 86 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=107090 $D=1
M487 477 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=111720 $D=1
M488 4 87 478 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=107090 $D=1
M489 8 87 479 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=111720 $D=1
M490 480 88 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=107090 $D=1
M491 481 88 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=111720 $D=1
M492 482 87 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=107090 $D=1
M493 483 87 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=111720 $D=1
M494 4 482 753 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=107090 $D=1
M495 8 483 754 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=111720 $D=1
M496 484 753 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=107090 $D=1
M497 485 754 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=111720 $D=1
M498 482 478 484 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=107090 $D=1
M499 483 479 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=111720 $D=1
M500 484 88 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=107090 $D=1
M501 485 88 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=111720 $D=1
M502 246 89 484 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=107090 $D=1
M503 247 89 485 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=111720 $D=1
M504 486 89 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=107090 $D=1
M505 487 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=111720 $D=1
M506 4 90 488 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=107090 $D=1
M507 8 90 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=111720 $D=1
M508 490 91 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=107090 $D=1
M509 491 91 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=111720 $D=1
M510 492 90 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=107090 $D=1
M511 493 90 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=111720 $D=1
M512 4 492 755 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=107090 $D=1
M513 8 493 756 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=111720 $D=1
M514 494 755 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=107090 $D=1
M515 495 756 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=111720 $D=1
M516 492 488 494 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=107090 $D=1
M517 493 489 495 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=111720 $D=1
M518 494 91 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=107090 $D=1
M519 495 91 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=111720 $D=1
M520 246 92 494 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=107090 $D=1
M521 247 92 495 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=111720 $D=1
M522 496 92 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=107090 $D=1
M523 497 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=111720 $D=1
M524 4 93 498 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=107090 $D=1
M525 8 93 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=111720 $D=1
M526 500 94 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=107090 $D=1
M527 501 94 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=111720 $D=1
M528 502 93 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=107090 $D=1
M529 503 93 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=111720 $D=1
M530 4 502 757 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=107090 $D=1
M531 8 503 758 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=111720 $D=1
M532 504 757 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=107090 $D=1
M533 505 758 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=111720 $D=1
M534 502 498 504 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=107090 $D=1
M535 503 499 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=111720 $D=1
M536 504 94 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=107090 $D=1
M537 505 94 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=111720 $D=1
M538 246 95 504 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=107090 $D=1
M539 247 95 505 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=111720 $D=1
M540 506 95 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=107090 $D=1
M541 507 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=111720 $D=1
M542 4 96 508 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=107090 $D=1
M543 8 96 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=111720 $D=1
M544 510 97 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=107090 $D=1
M545 511 97 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=111720 $D=1
M546 512 96 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=107090 $D=1
M547 513 96 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=111720 $D=1
M548 4 512 759 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=107090 $D=1
M549 8 513 760 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=111720 $D=1
M550 514 759 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=107090 $D=1
M551 515 760 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=111720 $D=1
M552 512 508 514 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=107090 $D=1
M553 513 509 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=111720 $D=1
M554 514 97 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=107090 $D=1
M555 515 97 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=111720 $D=1
M556 246 98 514 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=107090 $D=1
M557 247 98 515 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=111720 $D=1
M558 516 98 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=107090 $D=1
M559 517 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=111720 $D=1
M560 4 99 518 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=107090 $D=1
M561 8 99 519 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=111720 $D=1
M562 520 100 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=107090 $D=1
M563 521 100 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=111720 $D=1
M564 522 99 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=107090 $D=1
M565 523 99 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=111720 $D=1
M566 4 522 761 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=107090 $D=1
M567 8 523 762 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=111720 $D=1
M568 524 761 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=107090 $D=1
M569 525 762 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=111720 $D=1
M570 522 518 524 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=107090 $D=1
M571 523 519 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=111720 $D=1
M572 524 100 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=107090 $D=1
M573 525 100 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=111720 $D=1
M574 246 101 524 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=107090 $D=1
M575 247 101 525 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=111720 $D=1
M576 526 101 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=107090 $D=1
M577 527 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=111720 $D=1
M578 4 102 528 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=107090 $D=1
M579 8 102 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=111720 $D=1
M580 530 103 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=107090 $D=1
M581 531 103 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=111720 $D=1
M582 532 102 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=107090 $D=1
M583 533 102 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=111720 $D=1
M584 4 532 763 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=107090 $D=1
M585 8 533 764 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=111720 $D=1
M586 534 763 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=107090 $D=1
M587 535 764 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=111720 $D=1
M588 532 528 534 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=107090 $D=1
M589 533 529 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=111720 $D=1
M590 534 103 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=107090 $D=1
M591 535 103 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=111720 $D=1
M592 246 104 534 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=107090 $D=1
M593 247 104 535 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=111720 $D=1
M594 536 104 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=107090 $D=1
M595 537 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=111720 $D=1
M596 4 105 538 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=107090 $D=1
M597 8 105 539 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=111720 $D=1
M598 540 106 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=107090 $D=1
M599 541 106 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=111720 $D=1
M600 542 105 232 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=107090 $D=1
M601 543 105 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=111720 $D=1
M602 4 542 765 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=107090 $D=1
M603 8 543 766 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=111720 $D=1
M604 544 765 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=107090 $D=1
M605 545 766 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=111720 $D=1
M606 542 538 544 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=107090 $D=1
M607 543 539 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=111720 $D=1
M608 544 106 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=107090 $D=1
M609 545 106 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=111720 $D=1
M610 246 107 544 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=107090 $D=1
M611 247 107 545 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=111720 $D=1
M612 546 107 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=107090 $D=1
M613 547 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=111720 $D=1
M614 4 108 548 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=107090 $D=1
M615 8 108 549 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=111720 $D=1
M616 550 109 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=107090 $D=1
M617 551 109 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=111720 $D=1
M618 4 109 242 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=107090 $D=1
M619 8 109 243 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=111720 $D=1
M620 246 108 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=107090 $D=1
M621 247 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=111720 $D=1
M622 4 554 552 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=107090 $D=1
M623 8 555 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=111720 $D=1
M624 554 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=107090 $D=1
M625 555 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=111720 $D=1
M626 767 242 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=107090 $D=1
M627 768 243 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=111720 $D=1
M628 556 552 767 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=107090 $D=1
M629 557 553 768 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=111720 $D=1
M630 4 556 558 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=107090 $D=1
M631 8 557 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=111720 $D=1
M632 769 558 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=107090 $D=1
M633 770 559 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=111720 $D=1
M634 556 554 769 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=107090 $D=1
M635 557 555 770 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=111720 $D=1
M636 4 562 560 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=107090 $D=1
M637 8 563 561 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=111720 $D=1
M638 562 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=107090 $D=1
M639 563 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=111720 $D=1
M640 771 246 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=107090 $D=1
M641 772 247 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=111720 $D=1
M642 564 560 771 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=107090 $D=1
M643 565 561 772 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=111720 $D=1
M644 4 564 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=107090 $D=1
M645 8 565 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=111720 $D=1
M646 773 111 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=107090 $D=1
M647 774 112 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=111720 $D=1
M648 564 562 773 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=107090 $D=1
M649 565 563 774 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=111720 $D=1
M650 566 113 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=107090 $D=1
M651 567 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=111720 $D=1
M652 568 566 558 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=107090 $D=1
M653 569 567 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=111720 $D=1
M654 114 113 568 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=107090 $D=1
M655 114 113 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=111720 $D=1
M656 570 115 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=107090 $D=1
M657 571 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=111720 $D=1
M658 572 570 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=107090 $D=1
M659 573 571 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=111720 $D=1
M660 775 115 572 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=107090 $D=1
M661 776 115 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=111720 $D=1
M662 4 111 775 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=107090 $D=1
M663 8 112 776 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=111720 $D=1
M664 574 117 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=107090 $D=1
M665 575 117 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=111720 $D=1
M666 576 574 572 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=107090 $D=1
M667 577 575 573 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=111720 $D=1
M668 9 117 576 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=107090 $D=1
M669 10 117 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=111720 $D=1
M670 579 578 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=107090 $D=1
M671 580 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=111720 $D=1
M672 4 583 581 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=107090 $D=1
M673 8 584 582 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=111720 $D=1
M674 585 568 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=107090 $D=1
M675 586 569 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=111720 $D=1
M676 583 585 578 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=107090 $D=1
M677 584 586 119 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=111720 $D=1
M678 579 568 583 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=107090 $D=1
M679 580 569 584 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=111720 $D=1
M680 587 581 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=107090 $D=1
M681 588 582 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=111720 $D=1
M682 589 587 576 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=107090 $D=1
M683 578 588 577 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=111720 $D=1
M684 568 581 589 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=107090 $D=1
M685 569 582 578 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=111720 $D=1
M686 590 589 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=107090 $D=1
M687 591 578 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=111720 $D=1
M688 592 581 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=107090 $D=1
M689 593 582 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=111720 $D=1
M690 594 592 590 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=107090 $D=1
M691 595 593 591 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=111720 $D=1
M692 576 581 594 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=107090 $D=1
M693 577 582 595 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=111720 $D=1
M694 596 568 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=107090 $D=1
M695 597 569 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=111720 $D=1
M696 4 576 596 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=107090 $D=1
M697 8 577 597 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=111720 $D=1
M698 598 594 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=107090 $D=1
M699 599 595 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=111720 $D=1
M700 795 568 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=107090 $D=1
M701 796 569 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=111720 $D=1
M702 600 576 795 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=107090 $D=1
M703 601 577 796 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=111720 $D=1
M704 797 568 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=107090 $D=1
M705 798 569 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=111720 $D=1
M706 602 576 797 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=107090 $D=1
M707 603 577 798 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=111720 $D=1
M708 606 568 604 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=107090 $D=1
M709 607 569 605 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=111720 $D=1
M710 604 576 606 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=107090 $D=1
M711 605 577 607 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=111720 $D=1
M712 4 602 604 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=107090 $D=1
M713 8 603 605 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=111720 $D=1
M714 608 124 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=107090 $D=1
M715 609 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=111720 $D=1
M716 610 608 596 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=107090 $D=1
M717 611 609 597 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=111720 $D=1
M718 600 124 610 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=107090 $D=1
M719 601 124 611 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=111720 $D=1
M720 612 608 598 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=107090 $D=1
M721 613 609 599 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=111720 $D=1
M722 606 124 612 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=107090 $D=1
M723 607 124 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=111720 $D=1
M724 614 125 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=107090 $D=1
M725 615 125 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=111720 $D=1
M726 616 614 612 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=107090 $D=1
M727 617 615 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=111720 $D=1
M728 610 125 616 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=107090 $D=1
M729 611 125 617 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=111720 $D=1
M730 11 616 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=107090 $D=1
M731 12 617 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=111720 $D=1
M732 618 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=107090 $D=1
M733 619 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=111720 $D=1
M734 620 618 127 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=107090 $D=1
M735 621 619 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=111720 $D=1
M736 129 126 620 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=107090 $D=1
M737 130 126 621 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=111720 $D=1
M738 622 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=107090 $D=1
M739 623 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=111720 $D=1
M740 624 622 131 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=107090 $D=1
M741 625 623 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=111720 $D=1
M742 133 126 624 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=107090 $D=1
M743 134 126 625 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=111720 $D=1
M744 626 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=107090 $D=1
M745 627 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=111720 $D=1
M746 137 626 135 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=107090 $D=1
M747 137 627 136 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=111720 $D=1
M748 116 126 137 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=107090 $D=1
M749 122 126 137 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=111720 $D=1
M750 628 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=107090 $D=1
M751 629 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=111720 $D=1
M752 630 628 138 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=107090 $D=1
M753 631 629 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=111720 $D=1
M754 118 126 630 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=107090 $D=1
M755 139 126 631 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=111720 $D=1
M756 632 126 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=107090 $D=1
M757 633 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=111720 $D=1
M758 634 632 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=107090 $D=1
M759 635 633 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=111720 $D=1
M760 140 126 634 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=107090 $D=1
M761 141 126 635 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=111720 $D=1
M762 4 568 777 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=107090 $D=1
M763 8 569 778 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=111720 $D=1
M764 130 777 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=107090 $D=1
M765 127 778 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=111720 $D=1
M766 636 142 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=107090 $D=1
M767 637 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=111720 $D=1
M768 143 636 130 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=107090 $D=1
M769 144 637 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=111720 $D=1
M770 620 142 143 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=107090 $D=1
M771 621 142 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=111720 $D=1
M772 638 145 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=107090 $D=1
M773 639 145 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=111720 $D=1
M774 123 638 143 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=107090 $D=1
M775 146 639 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=111720 $D=1
M776 624 145 123 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=107090 $D=1
M777 625 145 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=111720 $D=1
M778 640 147 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=107090 $D=1
M779 641 147 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=111720 $D=1
M780 120 640 123 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=107090 $D=1
M781 121 641 146 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=111720 $D=1
M782 137 147 120 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=107090 $D=1
M783 137 147 121 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=111720 $D=1
M784 642 148 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=107090 $D=1
M785 643 148 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=111720 $D=1
M786 149 642 120 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=107090 $D=1
M787 150 643 121 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=111720 $D=1
M788 630 148 149 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=107090 $D=1
M789 631 148 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=111720 $D=1
M790 644 151 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=107090 $D=1
M791 645 151 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=111720 $D=1
M792 218 644 149 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=107090 $D=1
M793 219 645 150 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=111720 $D=1
M794 634 151 218 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=107090 $D=1
M795 635 151 219 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=111720 $D=1
M796 646 152 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=107090 $D=1
M797 647 152 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=111720 $D=1
M798 648 646 111 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=107090 $D=1
M799 649 647 112 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=111720 $D=1
M800 9 152 648 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=107090 $D=1
M801 10 152 649 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=111720 $D=1
M802 799 558 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=107090 $D=1
M803 800 559 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=111720 $D=1
M804 650 648 799 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=107090 $D=1
M805 651 649 800 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=111720 $D=1
M806 654 558 652 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=107090 $D=1
M807 655 559 653 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=111720 $D=1
M808 652 648 654 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=107090 $D=1
M809 653 649 655 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=111720 $D=1
M810 4 650 652 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=107090 $D=1
M811 8 651 653 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=111720 $D=1
M812 801 153 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=107090 $D=1
M813 802 656 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=111720 $D=1
M814 779 654 801 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=107090 $D=1
M815 780 655 802 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=111720 $D=1
M816 656 779 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=107090 $D=1
M817 154 780 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=111720 $D=1
M818 657 558 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=107090 $D=1
M819 658 559 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=111720 $D=1
M820 4 659 657 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=107090 $D=1
M821 8 660 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=111720 $D=1
M822 659 648 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=107090 $D=1
M823 660 649 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=111720 $D=1
M824 803 657 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=107090 $D=1
M825 804 658 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=111720 $D=1
M826 661 153 803 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=107090 $D=1
M827 662 656 804 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=111720 $D=1
M828 664 155 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=107090 $D=1
M829 665 663 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=111720 $D=1
M830 805 661 4 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=107090 $D=1
M831 806 662 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=111720 $D=1
M832 663 664 805 4 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=107090 $D=1
M833 156 665 806 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=111720 $D=1
M834 667 666 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=107090 $D=1
M835 668 157 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=111720 $D=1
M836 4 671 669 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=107090 $D=1
M837 8 672 670 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=111720 $D=1
M838 673 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=107090 $D=1
M839 674 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=111720 $D=1
M840 671 673 666 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=107090 $D=1
M841 672 674 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=111720 $D=1
M842 667 114 671 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=107090 $D=1
M843 668 114 672 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=111720 $D=1
M844 675 669 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=107090 $D=1
M845 676 670 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=111720 $D=1
M846 158 675 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=107090 $D=1
M847 666 676 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=111720 $D=1
M848 114 669 158 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=107090 $D=1
M849 114 670 666 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=111720 $D=1
M850 677 158 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=107090 $D=1
M851 678 666 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=111720 $D=1
M852 679 669 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=107090 $D=1
M853 680 670 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=111720 $D=1
M854 220 679 677 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=107090 $D=1
M855 221 680 678 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=111720 $D=1
M856 4 669 220 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=107090 $D=1
M857 8 670 221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=111720 $D=1
M858 681 159 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=107090 $D=1
M859 682 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=111720 $D=1
M860 683 681 220 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=107090 $D=1
M861 684 682 221 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=111720 $D=1
M862 11 159 683 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=107090 $D=1
M863 12 159 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=111720 $D=1
M864 685 160 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=107090 $D=1
M865 686 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=111720 $D=1
M866 160 685 683 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=107090 $D=1
M867 160 686 684 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=111720 $D=1
M868 4 160 160 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=107090 $D=1
M869 8 160 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=111720 $D=1
M870 687 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=107090 $D=1
M871 688 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=111720 $D=1
M872 4 687 689 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=107090 $D=1
M873 8 688 690 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=111720 $D=1
M874 691 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=107090 $D=1
M875 692 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=111720 $D=1
M876 693 687 160 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=107090 $D=1
M877 694 688 160 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=111720 $D=1
M878 4 693 781 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=107090 $D=1
M879 8 694 782 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=111720 $D=1
M880 695 781 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=107090 $D=1
M881 696 782 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=111720 $D=1
M882 693 689 695 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=107090 $D=1
M883 694 690 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=111720 $D=1
M884 697 110 695 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=107090 $D=1
M885 698 110 696 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=111720 $D=1
M886 4 701 699 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=107090 $D=1
M887 8 702 700 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=111720 $D=1
M888 701 110 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=107090 $D=1
M889 702 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=111720 $D=1
M890 783 697 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=107090 $D=1
M891 784 698 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=111720 $D=1
M892 703 699 783 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=107090 $D=1
M893 704 700 784 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=111720 $D=1
M894 4 703 114 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=107090 $D=1
M895 8 704 114 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=111720 $D=1
M896 785 114 4 4 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=107090 $D=1
M897 786 114 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=111720 $D=1
M898 703 701 785 4 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=107090 $D=1
M899 704 702 786 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=111720 $D=1
M900 194 1 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=108340 $D=0
M901 195 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=112970 $D=0
M902 196 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=108340 $D=0
M903 197 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=112970 $D=0
M904 4 194 196 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=108340 $D=0
M905 8 195 197 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=112970 $D=0
M906 198 1 3 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=108340 $D=0
M907 199 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=112970 $D=0
M908 2 194 198 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=108340 $D=0
M909 3 195 199 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=112970 $D=0
M910 200 1 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=108340 $D=0
M911 201 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=112970 $D=0
M912 2 194 200 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=108340 $D=0
M913 3 195 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=112970 $D=0
M914 204 5 200 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=108340 $D=0
M915 205 5 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=112970 $D=0
M916 202 5 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=108340 $D=0
M917 203 5 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=112970 $D=0
M918 206 5 198 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=108340 $D=0
M919 207 5 199 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=112970 $D=0
M920 196 202 206 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=108340 $D=0
M921 197 203 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=112970 $D=0
M922 208 6 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=108340 $D=0
M923 209 6 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=112970 $D=0
M924 210 6 206 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=108340 $D=0
M925 211 6 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=112970 $D=0
M926 204 208 210 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=108340 $D=0
M927 205 209 211 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=112970 $D=0
M928 212 7 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=108340 $D=0
M929 213 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=112970 $D=0
M930 214 7 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=108340 $D=0
M931 215 7 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=112970 $D=0
M932 9 212 214 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=108340 $D=0
M933 10 213 215 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=112970 $D=0
M934 216 7 11 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=108340 $D=0
M935 217 7 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=112970 $D=0
M936 218 212 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=108340 $D=0
M937 219 213 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=112970 $D=0
M938 222 7 220 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=108340 $D=0
M939 223 7 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=112970 $D=0
M940 210 212 222 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=108340 $D=0
M941 211 213 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=112970 $D=0
M942 226 13 222 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=108340 $D=0
M943 227 13 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=112970 $D=0
M944 224 13 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=108340 $D=0
M945 225 13 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=112970 $D=0
M946 228 13 216 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=108340 $D=0
M947 229 13 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=112970 $D=0
M948 214 224 228 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=108340 $D=0
M949 215 225 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=112970 $D=0
M950 230 14 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=108340 $D=0
M951 231 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=112970 $D=0
M952 232 14 228 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=108340 $D=0
M953 233 14 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=112970 $D=0
M954 226 230 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=108340 $D=0
M955 227 231 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=112970 $D=0
M956 161 15 234 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=108340 $D=0
M957 162 15 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=112970 $D=0
M958 236 16 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=108340 $D=0
M959 237 16 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=112970 $D=0
M960 238 234 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=108340 $D=0
M961 239 235 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=112970 $D=0
M962 161 238 705 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=108340 $D=0
M963 162 239 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=112970 $D=0
M964 240 705 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=108340 $D=0
M965 241 706 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=112970 $D=0
M966 238 15 240 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=108340 $D=0
M967 239 15 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=112970 $D=0
M968 240 236 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=108340 $D=0
M969 241 237 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=112970 $D=0
M970 246 244 240 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=108340 $D=0
M971 247 245 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=112970 $D=0
M972 244 17 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=108340 $D=0
M973 245 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=112970 $D=0
M974 161 18 248 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=108340 $D=0
M975 162 18 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=112970 $D=0
M976 250 19 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=108340 $D=0
M977 251 19 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=112970 $D=0
M978 252 248 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=108340 $D=0
M979 253 249 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=112970 $D=0
M980 161 252 707 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=108340 $D=0
M981 162 253 708 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=112970 $D=0
M982 254 707 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=108340 $D=0
M983 255 708 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=112970 $D=0
M984 252 18 254 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=108340 $D=0
M985 253 18 255 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=112970 $D=0
M986 254 250 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=108340 $D=0
M987 255 251 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=112970 $D=0
M988 246 256 254 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=108340 $D=0
M989 247 257 255 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=112970 $D=0
M990 256 20 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=108340 $D=0
M991 257 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=112970 $D=0
M992 161 21 258 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=108340 $D=0
M993 162 21 259 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=112970 $D=0
M994 260 22 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=108340 $D=0
M995 261 22 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=112970 $D=0
M996 262 258 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=108340 $D=0
M997 263 259 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=112970 $D=0
M998 161 262 709 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=108340 $D=0
M999 162 263 710 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=112970 $D=0
M1000 264 709 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=108340 $D=0
M1001 265 710 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=112970 $D=0
M1002 262 21 264 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=108340 $D=0
M1003 263 21 265 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=112970 $D=0
M1004 264 260 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=108340 $D=0
M1005 265 261 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=112970 $D=0
M1006 246 266 264 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=108340 $D=0
M1007 247 267 265 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=112970 $D=0
M1008 266 23 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=108340 $D=0
M1009 267 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=112970 $D=0
M1010 161 24 268 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=108340 $D=0
M1011 162 24 269 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=112970 $D=0
M1012 270 25 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=108340 $D=0
M1013 271 25 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=112970 $D=0
M1014 272 268 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=108340 $D=0
M1015 273 269 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=112970 $D=0
M1016 161 272 711 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=108340 $D=0
M1017 162 273 712 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=112970 $D=0
M1018 274 711 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=108340 $D=0
M1019 275 712 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=112970 $D=0
M1020 272 24 274 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=108340 $D=0
M1021 273 24 275 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=112970 $D=0
M1022 274 270 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=108340 $D=0
M1023 275 271 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=112970 $D=0
M1024 246 276 274 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=108340 $D=0
M1025 247 277 275 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=112970 $D=0
M1026 276 26 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=108340 $D=0
M1027 277 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=112970 $D=0
M1028 161 27 278 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=108340 $D=0
M1029 162 27 279 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=112970 $D=0
M1030 280 28 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=108340 $D=0
M1031 281 28 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=112970 $D=0
M1032 282 278 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=108340 $D=0
M1033 283 279 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=112970 $D=0
M1034 161 282 713 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=108340 $D=0
M1035 162 283 714 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=112970 $D=0
M1036 284 713 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=108340 $D=0
M1037 285 714 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=112970 $D=0
M1038 282 27 284 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=108340 $D=0
M1039 283 27 285 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=112970 $D=0
M1040 284 280 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=108340 $D=0
M1041 285 281 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=112970 $D=0
M1042 246 286 284 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=108340 $D=0
M1043 247 287 285 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=112970 $D=0
M1044 286 29 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=108340 $D=0
M1045 287 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=112970 $D=0
M1046 161 30 288 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=108340 $D=0
M1047 162 30 289 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=112970 $D=0
M1048 290 31 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=108340 $D=0
M1049 291 31 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=112970 $D=0
M1050 292 288 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=108340 $D=0
M1051 293 289 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=112970 $D=0
M1052 161 292 715 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=108340 $D=0
M1053 162 293 716 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=112970 $D=0
M1054 294 715 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=108340 $D=0
M1055 295 716 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=112970 $D=0
M1056 292 30 294 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=108340 $D=0
M1057 293 30 295 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=112970 $D=0
M1058 294 290 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=108340 $D=0
M1059 295 291 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=112970 $D=0
M1060 246 296 294 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=108340 $D=0
M1061 247 297 295 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=112970 $D=0
M1062 296 32 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=108340 $D=0
M1063 297 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=112970 $D=0
M1064 161 33 298 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=108340 $D=0
M1065 162 33 299 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=112970 $D=0
M1066 300 34 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=108340 $D=0
M1067 301 34 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=112970 $D=0
M1068 302 298 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=108340 $D=0
M1069 303 299 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=112970 $D=0
M1070 161 302 717 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=108340 $D=0
M1071 162 303 718 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=112970 $D=0
M1072 304 717 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=108340 $D=0
M1073 305 718 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=112970 $D=0
M1074 302 33 304 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=108340 $D=0
M1075 303 33 305 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=112970 $D=0
M1076 304 300 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=108340 $D=0
M1077 305 301 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=112970 $D=0
M1078 246 306 304 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=108340 $D=0
M1079 247 307 305 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=112970 $D=0
M1080 306 35 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=108340 $D=0
M1081 307 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=112970 $D=0
M1082 161 36 308 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=108340 $D=0
M1083 162 36 309 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=112970 $D=0
M1084 310 37 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=108340 $D=0
M1085 311 37 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=112970 $D=0
M1086 312 308 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=108340 $D=0
M1087 313 309 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=112970 $D=0
M1088 161 312 719 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=108340 $D=0
M1089 162 313 720 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=112970 $D=0
M1090 314 719 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=108340 $D=0
M1091 315 720 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=112970 $D=0
M1092 312 36 314 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=108340 $D=0
M1093 313 36 315 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=112970 $D=0
M1094 314 310 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=108340 $D=0
M1095 315 311 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=112970 $D=0
M1096 246 316 314 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=108340 $D=0
M1097 247 317 315 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=112970 $D=0
M1098 316 38 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=108340 $D=0
M1099 317 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=112970 $D=0
M1100 161 39 318 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=108340 $D=0
M1101 162 39 319 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=112970 $D=0
M1102 320 40 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=108340 $D=0
M1103 321 40 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=112970 $D=0
M1104 322 318 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=108340 $D=0
M1105 323 319 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=112970 $D=0
M1106 161 322 721 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=108340 $D=0
M1107 162 323 722 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=112970 $D=0
M1108 324 721 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=108340 $D=0
M1109 325 722 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=112970 $D=0
M1110 322 39 324 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=108340 $D=0
M1111 323 39 325 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=112970 $D=0
M1112 324 320 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=108340 $D=0
M1113 325 321 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=112970 $D=0
M1114 246 326 324 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=108340 $D=0
M1115 247 327 325 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=112970 $D=0
M1116 326 41 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=108340 $D=0
M1117 327 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=112970 $D=0
M1118 161 42 328 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=108340 $D=0
M1119 162 42 329 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=112970 $D=0
M1120 330 43 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=108340 $D=0
M1121 331 43 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=112970 $D=0
M1122 332 328 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=108340 $D=0
M1123 333 329 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=112970 $D=0
M1124 161 332 723 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=108340 $D=0
M1125 162 333 724 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=112970 $D=0
M1126 334 723 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=108340 $D=0
M1127 335 724 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=112970 $D=0
M1128 332 42 334 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=108340 $D=0
M1129 333 42 335 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=112970 $D=0
M1130 334 330 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=108340 $D=0
M1131 335 331 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=112970 $D=0
M1132 246 336 334 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=108340 $D=0
M1133 247 337 335 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=112970 $D=0
M1134 336 44 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=108340 $D=0
M1135 337 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=112970 $D=0
M1136 161 45 338 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=108340 $D=0
M1137 162 45 339 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=112970 $D=0
M1138 340 46 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=108340 $D=0
M1139 341 46 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=112970 $D=0
M1140 342 338 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=108340 $D=0
M1141 343 339 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=112970 $D=0
M1142 161 342 725 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=108340 $D=0
M1143 162 343 726 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=112970 $D=0
M1144 344 725 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=108340 $D=0
M1145 345 726 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=112970 $D=0
M1146 342 45 344 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=108340 $D=0
M1147 343 45 345 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=112970 $D=0
M1148 344 340 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=108340 $D=0
M1149 345 341 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=112970 $D=0
M1150 246 346 344 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=108340 $D=0
M1151 247 347 345 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=112970 $D=0
M1152 346 47 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=108340 $D=0
M1153 347 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=112970 $D=0
M1154 161 48 348 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=108340 $D=0
M1155 162 48 349 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=112970 $D=0
M1156 350 49 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=108340 $D=0
M1157 351 49 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=112970 $D=0
M1158 352 348 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=108340 $D=0
M1159 353 349 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=112970 $D=0
M1160 161 352 727 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=108340 $D=0
M1161 162 353 728 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=112970 $D=0
M1162 354 727 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=108340 $D=0
M1163 355 728 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=112970 $D=0
M1164 352 48 354 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=108340 $D=0
M1165 353 48 355 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=112970 $D=0
M1166 354 350 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=108340 $D=0
M1167 355 351 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=112970 $D=0
M1168 246 356 354 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=108340 $D=0
M1169 247 357 355 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=112970 $D=0
M1170 356 50 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=108340 $D=0
M1171 357 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=112970 $D=0
M1172 161 51 358 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=108340 $D=0
M1173 162 51 359 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=112970 $D=0
M1174 360 52 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=108340 $D=0
M1175 361 52 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=112970 $D=0
M1176 362 358 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=108340 $D=0
M1177 363 359 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=112970 $D=0
M1178 161 362 729 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=108340 $D=0
M1179 162 363 730 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=112970 $D=0
M1180 364 729 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=108340 $D=0
M1181 365 730 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=112970 $D=0
M1182 362 51 364 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=108340 $D=0
M1183 363 51 365 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=112970 $D=0
M1184 364 360 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=108340 $D=0
M1185 365 361 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=112970 $D=0
M1186 246 366 364 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=108340 $D=0
M1187 247 367 365 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=112970 $D=0
M1188 366 53 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=108340 $D=0
M1189 367 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=112970 $D=0
M1190 161 54 368 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=108340 $D=0
M1191 162 54 369 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=112970 $D=0
M1192 370 55 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=108340 $D=0
M1193 371 55 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=112970 $D=0
M1194 372 368 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=108340 $D=0
M1195 373 369 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=112970 $D=0
M1196 161 372 731 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=108340 $D=0
M1197 162 373 732 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=112970 $D=0
M1198 374 731 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=108340 $D=0
M1199 375 732 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=112970 $D=0
M1200 372 54 374 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=108340 $D=0
M1201 373 54 375 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=112970 $D=0
M1202 374 370 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=108340 $D=0
M1203 375 371 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=112970 $D=0
M1204 246 376 374 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=108340 $D=0
M1205 247 377 375 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=112970 $D=0
M1206 376 56 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=108340 $D=0
M1207 377 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=112970 $D=0
M1208 161 57 378 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=108340 $D=0
M1209 162 57 379 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=112970 $D=0
M1210 380 58 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=108340 $D=0
M1211 381 58 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=112970 $D=0
M1212 382 378 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=108340 $D=0
M1213 383 379 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=112970 $D=0
M1214 161 382 733 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=108340 $D=0
M1215 162 383 734 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=112970 $D=0
M1216 384 733 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=108340 $D=0
M1217 385 734 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=112970 $D=0
M1218 382 57 384 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=108340 $D=0
M1219 383 57 385 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=112970 $D=0
M1220 384 380 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=108340 $D=0
M1221 385 381 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=112970 $D=0
M1222 246 386 384 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=108340 $D=0
M1223 247 387 385 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=112970 $D=0
M1224 386 59 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=108340 $D=0
M1225 387 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=112970 $D=0
M1226 161 60 388 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=108340 $D=0
M1227 162 60 389 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=112970 $D=0
M1228 390 61 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=108340 $D=0
M1229 391 61 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=112970 $D=0
M1230 392 388 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=108340 $D=0
M1231 393 389 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=112970 $D=0
M1232 161 392 735 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=108340 $D=0
M1233 162 393 736 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=112970 $D=0
M1234 394 735 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=108340 $D=0
M1235 395 736 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=112970 $D=0
M1236 392 60 394 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=108340 $D=0
M1237 393 60 395 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=112970 $D=0
M1238 394 390 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=108340 $D=0
M1239 395 391 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=112970 $D=0
M1240 246 396 394 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=108340 $D=0
M1241 247 397 395 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=112970 $D=0
M1242 396 62 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=108340 $D=0
M1243 397 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=112970 $D=0
M1244 161 63 398 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=108340 $D=0
M1245 162 63 399 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=112970 $D=0
M1246 400 64 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=108340 $D=0
M1247 401 64 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=112970 $D=0
M1248 402 398 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=108340 $D=0
M1249 403 399 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=112970 $D=0
M1250 161 402 737 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=108340 $D=0
M1251 162 403 738 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=112970 $D=0
M1252 404 737 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=108340 $D=0
M1253 405 738 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=112970 $D=0
M1254 402 63 404 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=108340 $D=0
M1255 403 63 405 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=112970 $D=0
M1256 404 400 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=108340 $D=0
M1257 405 401 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=112970 $D=0
M1258 246 406 404 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=108340 $D=0
M1259 247 407 405 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=112970 $D=0
M1260 406 65 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=108340 $D=0
M1261 407 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=112970 $D=0
M1262 161 66 408 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=108340 $D=0
M1263 162 66 409 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=112970 $D=0
M1264 410 67 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=108340 $D=0
M1265 411 67 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=112970 $D=0
M1266 412 408 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=108340 $D=0
M1267 413 409 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=112970 $D=0
M1268 161 412 739 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=108340 $D=0
M1269 162 413 740 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=112970 $D=0
M1270 414 739 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=108340 $D=0
M1271 415 740 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=112970 $D=0
M1272 412 66 414 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=108340 $D=0
M1273 413 66 415 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=112970 $D=0
M1274 414 410 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=108340 $D=0
M1275 415 411 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=112970 $D=0
M1276 246 416 414 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=108340 $D=0
M1277 247 417 415 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=112970 $D=0
M1278 416 68 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=108340 $D=0
M1279 417 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=112970 $D=0
M1280 161 69 418 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=108340 $D=0
M1281 162 69 419 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=112970 $D=0
M1282 420 70 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=108340 $D=0
M1283 421 70 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=112970 $D=0
M1284 422 418 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=108340 $D=0
M1285 423 419 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=112970 $D=0
M1286 161 422 741 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=108340 $D=0
M1287 162 423 742 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=112970 $D=0
M1288 424 741 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=108340 $D=0
M1289 425 742 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=112970 $D=0
M1290 422 69 424 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=108340 $D=0
M1291 423 69 425 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=112970 $D=0
M1292 424 420 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=108340 $D=0
M1293 425 421 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=112970 $D=0
M1294 246 426 424 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=108340 $D=0
M1295 247 427 425 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=112970 $D=0
M1296 426 71 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=108340 $D=0
M1297 427 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=112970 $D=0
M1298 161 72 428 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=108340 $D=0
M1299 162 72 429 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=112970 $D=0
M1300 430 73 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=108340 $D=0
M1301 431 73 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=112970 $D=0
M1302 432 428 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=108340 $D=0
M1303 433 429 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=112970 $D=0
M1304 161 432 743 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=108340 $D=0
M1305 162 433 744 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=112970 $D=0
M1306 434 743 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=108340 $D=0
M1307 435 744 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=112970 $D=0
M1308 432 72 434 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=108340 $D=0
M1309 433 72 435 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=112970 $D=0
M1310 434 430 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=108340 $D=0
M1311 435 431 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=112970 $D=0
M1312 246 436 434 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=108340 $D=0
M1313 247 437 435 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=112970 $D=0
M1314 436 74 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=108340 $D=0
M1315 437 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=112970 $D=0
M1316 161 75 438 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=108340 $D=0
M1317 162 75 439 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=112970 $D=0
M1318 440 76 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=108340 $D=0
M1319 441 76 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=112970 $D=0
M1320 442 438 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=108340 $D=0
M1321 443 439 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=112970 $D=0
M1322 161 442 745 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=108340 $D=0
M1323 162 443 746 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=112970 $D=0
M1324 444 745 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=108340 $D=0
M1325 445 746 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=112970 $D=0
M1326 442 75 444 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=108340 $D=0
M1327 443 75 445 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=112970 $D=0
M1328 444 440 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=108340 $D=0
M1329 445 441 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=112970 $D=0
M1330 246 446 444 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=108340 $D=0
M1331 247 447 445 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=112970 $D=0
M1332 446 77 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=108340 $D=0
M1333 447 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=112970 $D=0
M1334 161 78 448 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=108340 $D=0
M1335 162 78 449 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=112970 $D=0
M1336 450 79 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=108340 $D=0
M1337 451 79 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=112970 $D=0
M1338 452 448 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=108340 $D=0
M1339 453 449 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=112970 $D=0
M1340 161 452 747 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=108340 $D=0
M1341 162 453 748 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=112970 $D=0
M1342 454 747 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=108340 $D=0
M1343 455 748 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=112970 $D=0
M1344 452 78 454 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=108340 $D=0
M1345 453 78 455 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=112970 $D=0
M1346 454 450 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=108340 $D=0
M1347 455 451 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=112970 $D=0
M1348 246 456 454 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=108340 $D=0
M1349 247 457 455 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=112970 $D=0
M1350 456 80 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=108340 $D=0
M1351 457 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=112970 $D=0
M1352 161 81 458 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=108340 $D=0
M1353 162 81 459 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=112970 $D=0
M1354 460 82 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=108340 $D=0
M1355 461 82 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=112970 $D=0
M1356 462 458 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=108340 $D=0
M1357 463 459 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=112970 $D=0
M1358 161 462 749 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=108340 $D=0
M1359 162 463 750 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=112970 $D=0
M1360 464 749 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=108340 $D=0
M1361 465 750 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=112970 $D=0
M1362 462 81 464 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=108340 $D=0
M1363 463 81 465 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=112970 $D=0
M1364 464 460 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=108340 $D=0
M1365 465 461 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=112970 $D=0
M1366 246 466 464 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=108340 $D=0
M1367 247 467 465 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=112970 $D=0
M1368 466 83 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=108340 $D=0
M1369 467 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=112970 $D=0
M1370 161 84 468 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=108340 $D=0
M1371 162 84 469 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=112970 $D=0
M1372 470 85 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=108340 $D=0
M1373 471 85 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=112970 $D=0
M1374 472 468 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=108340 $D=0
M1375 473 469 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=112970 $D=0
M1376 161 472 751 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=108340 $D=0
M1377 162 473 752 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=112970 $D=0
M1378 474 751 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=108340 $D=0
M1379 475 752 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=112970 $D=0
M1380 472 84 474 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=108340 $D=0
M1381 473 84 475 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=112970 $D=0
M1382 474 470 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=108340 $D=0
M1383 475 471 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=112970 $D=0
M1384 246 476 474 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=108340 $D=0
M1385 247 477 475 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=112970 $D=0
M1386 476 86 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=108340 $D=0
M1387 477 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=112970 $D=0
M1388 161 87 478 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=108340 $D=0
M1389 162 87 479 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=112970 $D=0
M1390 480 88 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=108340 $D=0
M1391 481 88 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=112970 $D=0
M1392 482 478 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=108340 $D=0
M1393 483 479 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=112970 $D=0
M1394 161 482 753 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=108340 $D=0
M1395 162 483 754 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=112970 $D=0
M1396 484 753 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=108340 $D=0
M1397 485 754 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=112970 $D=0
M1398 482 87 484 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=108340 $D=0
M1399 483 87 485 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=112970 $D=0
M1400 484 480 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=108340 $D=0
M1401 485 481 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=112970 $D=0
M1402 246 486 484 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=108340 $D=0
M1403 247 487 485 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=112970 $D=0
M1404 486 89 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=108340 $D=0
M1405 487 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=112970 $D=0
M1406 161 90 488 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=108340 $D=0
M1407 162 90 489 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=112970 $D=0
M1408 490 91 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=108340 $D=0
M1409 491 91 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=112970 $D=0
M1410 492 488 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=108340 $D=0
M1411 493 489 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=112970 $D=0
M1412 161 492 755 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=108340 $D=0
M1413 162 493 756 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=112970 $D=0
M1414 494 755 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=108340 $D=0
M1415 495 756 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=112970 $D=0
M1416 492 90 494 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=108340 $D=0
M1417 493 90 495 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=112970 $D=0
M1418 494 490 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=108340 $D=0
M1419 495 491 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=112970 $D=0
M1420 246 496 494 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=108340 $D=0
M1421 247 497 495 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=112970 $D=0
M1422 496 92 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=108340 $D=0
M1423 497 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=112970 $D=0
M1424 161 93 498 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=108340 $D=0
M1425 162 93 499 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=112970 $D=0
M1426 500 94 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=108340 $D=0
M1427 501 94 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=112970 $D=0
M1428 502 498 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=108340 $D=0
M1429 503 499 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=112970 $D=0
M1430 161 502 757 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=108340 $D=0
M1431 162 503 758 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=112970 $D=0
M1432 504 757 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=108340 $D=0
M1433 505 758 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=112970 $D=0
M1434 502 93 504 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=108340 $D=0
M1435 503 93 505 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=112970 $D=0
M1436 504 500 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=108340 $D=0
M1437 505 501 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=112970 $D=0
M1438 246 506 504 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=108340 $D=0
M1439 247 507 505 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=112970 $D=0
M1440 506 95 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=108340 $D=0
M1441 507 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=112970 $D=0
M1442 161 96 508 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=108340 $D=0
M1443 162 96 509 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=112970 $D=0
M1444 510 97 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=108340 $D=0
M1445 511 97 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=112970 $D=0
M1446 512 508 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=108340 $D=0
M1447 513 509 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=112970 $D=0
M1448 161 512 759 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=108340 $D=0
M1449 162 513 760 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=112970 $D=0
M1450 514 759 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=108340 $D=0
M1451 515 760 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=112970 $D=0
M1452 512 96 514 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=108340 $D=0
M1453 513 96 515 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=112970 $D=0
M1454 514 510 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=108340 $D=0
M1455 515 511 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=112970 $D=0
M1456 246 516 514 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=108340 $D=0
M1457 247 517 515 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=112970 $D=0
M1458 516 98 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=108340 $D=0
M1459 517 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=112970 $D=0
M1460 161 99 518 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=108340 $D=0
M1461 162 99 519 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=112970 $D=0
M1462 520 100 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=108340 $D=0
M1463 521 100 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=112970 $D=0
M1464 522 518 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=108340 $D=0
M1465 523 519 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=112970 $D=0
M1466 161 522 761 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=108340 $D=0
M1467 162 523 762 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=112970 $D=0
M1468 524 761 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=108340 $D=0
M1469 525 762 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=112970 $D=0
M1470 522 99 524 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=108340 $D=0
M1471 523 99 525 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=112970 $D=0
M1472 524 520 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=108340 $D=0
M1473 525 521 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=112970 $D=0
M1474 246 526 524 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=108340 $D=0
M1475 247 527 525 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=112970 $D=0
M1476 526 101 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=108340 $D=0
M1477 527 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=112970 $D=0
M1478 161 102 528 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=108340 $D=0
M1479 162 102 529 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=112970 $D=0
M1480 530 103 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=108340 $D=0
M1481 531 103 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=112970 $D=0
M1482 532 528 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=108340 $D=0
M1483 533 529 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=112970 $D=0
M1484 161 532 763 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=108340 $D=0
M1485 162 533 764 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=112970 $D=0
M1486 534 763 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=108340 $D=0
M1487 535 764 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=112970 $D=0
M1488 532 102 534 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=108340 $D=0
M1489 533 102 535 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=112970 $D=0
M1490 534 530 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=108340 $D=0
M1491 535 531 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=112970 $D=0
M1492 246 536 534 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=108340 $D=0
M1493 247 537 535 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=112970 $D=0
M1494 536 104 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=108340 $D=0
M1495 537 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=112970 $D=0
M1496 161 105 538 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=108340 $D=0
M1497 162 105 539 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=112970 $D=0
M1498 540 106 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=108340 $D=0
M1499 541 106 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=112970 $D=0
M1500 542 538 232 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=108340 $D=0
M1501 543 539 233 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=112970 $D=0
M1502 161 542 765 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=108340 $D=0
M1503 162 543 766 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=112970 $D=0
M1504 544 765 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=108340 $D=0
M1505 545 766 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=112970 $D=0
M1506 542 105 544 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=108340 $D=0
M1507 543 105 545 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=112970 $D=0
M1508 544 540 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=108340 $D=0
M1509 545 541 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=112970 $D=0
M1510 246 546 544 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=108340 $D=0
M1511 247 547 545 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=112970 $D=0
M1512 546 107 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=108340 $D=0
M1513 547 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=112970 $D=0
M1514 161 108 548 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=108340 $D=0
M1515 162 108 549 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=112970 $D=0
M1516 550 109 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=108340 $D=0
M1517 551 109 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=112970 $D=0
M1518 4 550 242 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=108340 $D=0
M1519 8 551 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=112970 $D=0
M1520 246 548 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=108340 $D=0
M1521 247 549 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=112970 $D=0
M1522 161 554 552 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=108340 $D=0
M1523 162 555 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=112970 $D=0
M1524 554 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=108340 $D=0
M1525 555 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=112970 $D=0
M1526 767 242 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=108340 $D=0
M1527 768 243 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=112970 $D=0
M1528 556 554 767 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=108340 $D=0
M1529 557 555 768 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=112970 $D=0
M1530 161 556 558 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=108340 $D=0
M1531 162 557 559 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=112970 $D=0
M1532 769 558 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=108340 $D=0
M1533 770 559 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=112970 $D=0
M1534 556 552 769 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=108340 $D=0
M1535 557 553 770 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=112970 $D=0
M1536 161 562 560 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=108340 $D=0
M1537 162 563 561 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=112970 $D=0
M1538 562 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=108340 $D=0
M1539 563 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=112970 $D=0
M1540 771 246 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=108340 $D=0
M1541 772 247 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=112970 $D=0
M1542 564 562 771 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=108340 $D=0
M1543 565 563 772 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=112970 $D=0
M1544 161 564 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=108340 $D=0
M1545 162 565 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=112970 $D=0
M1546 773 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=108340 $D=0
M1547 774 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=112970 $D=0
M1548 564 560 773 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=108340 $D=0
M1549 565 561 774 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=112970 $D=0
M1550 566 113 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=108340 $D=0
M1551 567 113 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=112970 $D=0
M1552 568 113 558 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=108340 $D=0
M1553 569 113 559 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=112970 $D=0
M1554 114 566 568 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=108340 $D=0
M1555 114 567 569 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=112970 $D=0
M1556 570 115 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=108340 $D=0
M1557 571 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=112970 $D=0
M1558 572 115 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=108340 $D=0
M1559 573 115 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=112970 $D=0
M1560 775 570 572 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=108340 $D=0
M1561 776 571 573 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=112970 $D=0
M1562 161 111 775 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=108340 $D=0
M1563 162 112 776 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=112970 $D=0
M1564 574 117 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=108340 $D=0
M1565 575 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=112970 $D=0
M1566 576 117 572 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=108340 $D=0
M1567 577 117 573 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=112970 $D=0
M1568 9 574 576 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=108340 $D=0
M1569 10 575 577 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=112970 $D=0
M1570 579 578 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=108340 $D=0
M1571 580 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=112970 $D=0
M1572 161 583 581 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=108340 $D=0
M1573 162 584 582 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=112970 $D=0
M1574 585 568 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=108340 $D=0
M1575 586 569 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=112970 $D=0
M1576 583 568 578 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=108340 $D=0
M1577 584 569 119 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=112970 $D=0
M1578 579 585 583 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=108340 $D=0
M1579 580 586 584 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=112970 $D=0
M1580 587 581 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=108340 $D=0
M1581 588 582 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=112970 $D=0
M1582 589 581 576 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=108340 $D=0
M1583 578 582 577 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=112970 $D=0
M1584 568 587 589 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=108340 $D=0
M1585 569 588 578 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=112970 $D=0
M1586 590 589 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=108340 $D=0
M1587 591 578 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=112970 $D=0
M1588 592 581 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=108340 $D=0
M1589 593 582 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=112970 $D=0
M1590 594 581 590 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=108340 $D=0
M1591 595 582 591 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=112970 $D=0
M1592 576 592 594 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=108340 $D=0
M1593 577 593 595 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=112970 $D=0
M1594 787 568 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=107980 $D=0
M1595 788 569 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=112610 $D=0
M1596 596 576 787 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=107980 $D=0
M1597 597 577 788 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=112610 $D=0
M1598 598 594 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=108340 $D=0
M1599 599 595 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=112970 $D=0
M1600 600 568 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=108340 $D=0
M1601 601 569 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=112970 $D=0
M1602 161 576 600 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=108340 $D=0
M1603 162 577 601 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=112970 $D=0
M1604 602 568 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=108340 $D=0
M1605 603 569 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=112970 $D=0
M1606 161 576 602 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=108340 $D=0
M1607 162 577 603 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=112970 $D=0
M1608 789 568 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=108160 $D=0
M1609 790 569 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=112790 $D=0
M1610 606 576 789 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=108160 $D=0
M1611 607 577 790 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=112790 $D=0
M1612 161 602 606 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=108340 $D=0
M1613 162 603 607 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=112970 $D=0
M1614 608 124 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=108340 $D=0
M1615 609 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=112970 $D=0
M1616 610 124 596 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=108340 $D=0
M1617 611 124 597 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=112970 $D=0
M1618 600 608 610 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=108340 $D=0
M1619 601 609 611 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=112970 $D=0
M1620 612 124 598 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=108340 $D=0
M1621 613 124 599 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=112970 $D=0
M1622 606 608 612 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=108340 $D=0
M1623 607 609 613 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=112970 $D=0
M1624 614 125 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=108340 $D=0
M1625 615 125 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=112970 $D=0
M1626 616 125 612 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=108340 $D=0
M1627 617 125 613 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=112970 $D=0
M1628 610 614 616 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=108340 $D=0
M1629 611 615 617 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=112970 $D=0
M1630 11 616 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=108340 $D=0
M1631 12 617 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=112970 $D=0
M1632 618 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=108340 $D=0
M1633 619 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=112970 $D=0
M1634 620 126 127 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=108340 $D=0
M1635 621 126 128 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=112970 $D=0
M1636 129 618 620 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=108340 $D=0
M1637 130 619 621 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=112970 $D=0
M1638 622 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=108340 $D=0
M1639 623 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=112970 $D=0
M1640 624 126 131 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=108340 $D=0
M1641 625 126 132 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=112970 $D=0
M1642 133 622 624 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=108340 $D=0
M1643 134 623 625 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=112970 $D=0
M1644 626 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=108340 $D=0
M1645 627 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=112970 $D=0
M1646 137 126 135 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=108340 $D=0
M1647 137 126 136 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=112970 $D=0
M1648 116 626 137 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=108340 $D=0
M1649 122 627 137 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=112970 $D=0
M1650 628 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=108340 $D=0
M1651 629 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=112970 $D=0
M1652 630 126 138 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=108340 $D=0
M1653 631 126 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=112970 $D=0
M1654 118 628 630 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=108340 $D=0
M1655 139 629 631 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=112970 $D=0
M1656 632 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=108340 $D=0
M1657 633 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=112970 $D=0
M1658 634 126 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=108340 $D=0
M1659 635 126 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=112970 $D=0
M1660 140 632 634 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=108340 $D=0
M1661 141 633 635 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=112970 $D=0
M1662 161 568 777 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=108340 $D=0
M1663 162 569 778 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=112970 $D=0
M1664 130 777 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=108340 $D=0
M1665 127 778 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=112970 $D=0
M1666 636 142 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=108340 $D=0
M1667 637 142 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=112970 $D=0
M1668 143 142 130 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=108340 $D=0
M1669 144 142 127 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=112970 $D=0
M1670 620 636 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=108340 $D=0
M1671 621 637 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=112970 $D=0
M1672 638 145 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=108340 $D=0
M1673 639 145 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=112970 $D=0
M1674 123 145 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=108340 $D=0
M1675 146 145 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=112970 $D=0
M1676 624 638 123 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=108340 $D=0
M1677 625 639 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=112970 $D=0
M1678 640 147 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=108340 $D=0
M1679 641 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=112970 $D=0
M1680 120 147 123 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=108340 $D=0
M1681 121 147 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=112970 $D=0
M1682 137 640 120 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=108340 $D=0
M1683 137 641 121 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=112970 $D=0
M1684 642 148 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=108340 $D=0
M1685 643 148 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=112970 $D=0
M1686 149 148 120 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=108340 $D=0
M1687 150 148 121 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=112970 $D=0
M1688 630 642 149 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=108340 $D=0
M1689 631 643 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=112970 $D=0
M1690 644 151 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=108340 $D=0
M1691 645 151 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=112970 $D=0
M1692 218 151 149 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=108340 $D=0
M1693 219 151 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=112970 $D=0
M1694 634 644 218 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=108340 $D=0
M1695 635 645 219 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=112970 $D=0
M1696 646 152 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=108340 $D=0
M1697 647 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=112970 $D=0
M1698 648 152 111 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=108340 $D=0
M1699 649 152 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=112970 $D=0
M1700 9 646 648 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=108340 $D=0
M1701 10 647 649 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=112970 $D=0
M1702 650 558 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=108340 $D=0
M1703 651 559 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=112970 $D=0
M1704 161 648 650 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=108340 $D=0
M1705 162 649 651 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=112970 $D=0
M1706 791 558 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=108160 $D=0
M1707 792 559 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=112790 $D=0
M1708 654 648 791 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=108160 $D=0
M1709 655 649 792 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=112790 $D=0
M1710 161 650 654 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=108340 $D=0
M1711 162 651 655 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=112970 $D=0
M1712 779 153 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=108340 $D=0
M1713 780 656 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=112970 $D=0
M1714 161 654 779 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=108340 $D=0
M1715 162 655 780 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=112970 $D=0
M1716 656 779 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=108340 $D=0
M1717 154 780 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=112970 $D=0
M1718 793 558 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=107980 $D=0
M1719 794 559 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=112610 $D=0
M1720 657 659 793 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=107980 $D=0
M1721 658 660 794 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=112610 $D=0
M1722 659 648 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=108340 $D=0
M1723 660 649 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=112970 $D=0
M1724 661 657 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=108340 $D=0
M1725 662 658 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=112970 $D=0
M1726 161 153 661 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=108340 $D=0
M1727 162 656 662 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=112970 $D=0
M1728 664 155 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=108340 $D=0
M1729 665 663 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=112970 $D=0
M1730 663 661 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=108340 $D=0
M1731 156 662 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=112970 $D=0
M1732 161 664 663 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=108340 $D=0
M1733 162 665 156 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=112970 $D=0
M1734 667 666 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=108340 $D=0
M1735 668 157 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=112970 $D=0
M1736 161 671 669 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=108340 $D=0
M1737 162 672 670 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=112970 $D=0
M1738 673 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=108340 $D=0
M1739 674 114 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=112970 $D=0
M1740 671 114 666 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=108340 $D=0
M1741 672 114 157 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=112970 $D=0
M1742 667 673 671 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=108340 $D=0
M1743 668 674 672 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=112970 $D=0
M1744 675 669 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=108340 $D=0
M1745 676 670 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=112970 $D=0
M1746 158 669 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=108340 $D=0
M1747 666 670 8 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=112970 $D=0
M1748 114 675 158 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=108340 $D=0
M1749 114 676 666 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=112970 $D=0
M1750 677 158 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=108340 $D=0
M1751 678 666 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=112970 $D=0
M1752 679 669 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=108340 $D=0
M1753 680 670 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=112970 $D=0
M1754 220 669 677 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=108340 $D=0
M1755 221 670 678 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=112970 $D=0
M1756 4 679 220 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=108340 $D=0
M1757 8 680 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=112970 $D=0
M1758 681 159 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=108340 $D=0
M1759 682 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=112970 $D=0
M1760 683 159 220 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=108340 $D=0
M1761 684 159 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=112970 $D=0
M1762 11 681 683 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=108340 $D=0
M1763 12 682 684 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=112970 $D=0
M1764 685 160 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=108340 $D=0
M1765 686 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=112970 $D=0
M1766 160 160 683 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=108340 $D=0
M1767 160 160 684 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=112970 $D=0
M1768 4 685 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=108340 $D=0
M1769 8 686 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=112970 $D=0
M1770 687 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=108340 $D=0
M1771 688 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=112970 $D=0
M1772 161 687 689 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=108340 $D=0
M1773 162 688 690 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=112970 $D=0
M1774 691 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=108340 $D=0
M1775 692 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=112970 $D=0
M1776 693 689 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=108340 $D=0
M1777 694 690 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=112970 $D=0
M1778 161 693 781 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=108340 $D=0
M1779 162 694 782 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=112970 $D=0
M1780 695 781 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=108340 $D=0
M1781 696 782 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=112970 $D=0
M1782 693 687 695 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=108340 $D=0
M1783 694 688 696 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=112970 $D=0
M1784 697 691 695 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=108340 $D=0
M1785 698 692 696 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=112970 $D=0
M1786 161 701 699 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=108340 $D=0
M1787 162 702 700 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=112970 $D=0
M1788 701 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=108340 $D=0
M1789 702 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=112970 $D=0
M1790 783 697 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=108340 $D=0
M1791 784 698 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=112970 $D=0
M1792 703 701 783 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=108340 $D=0
M1793 704 702 784 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=112970 $D=0
M1794 161 703 114 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=108340 $D=0
M1795 162 704 114 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=112970 $D=0
M1796 785 114 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=108340 $D=0
M1797 786 114 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=112970 $D=0
M1798 703 699 785 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=108340 $D=0
M1799 704 700 786 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=112970 $D=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=808 EP=163 IP=1514 FDC=1800
M0 197 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=97830 $D=1
M1 198 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=102460 $D=1
M2 199 197 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=97830 $D=1
M3 200 198 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=102460 $D=1
M4 5 1 199 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=97830 $D=1
M5 6 1 200 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=102460 $D=1
M6 201 197 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=97830 $D=1
M7 202 198 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=102460 $D=1
M8 2 1 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=97830 $D=1
M9 3 1 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=102460 $D=1
M10 203 197 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=97830 $D=1
M11 204 198 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=102460 $D=1
M12 2 1 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=97830 $D=1
M13 3 1 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=102460 $D=1
M14 207 205 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=97830 $D=1
M15 208 206 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=102460 $D=1
M16 205 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=97830 $D=1
M17 206 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=102460 $D=1
M18 209 205 201 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=97830 $D=1
M19 210 206 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=102460 $D=1
M20 199 7 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=97830 $D=1
M21 200 7 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=102460 $D=1
M22 211 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=97830 $D=1
M23 212 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=102460 $D=1
M24 213 211 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=97830 $D=1
M25 214 212 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=102460 $D=1
M26 207 8 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=97830 $D=1
M27 208 8 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=102460 $D=1
M28 215 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=97830 $D=1
M29 216 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=102460 $D=1
M30 217 215 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=97830 $D=1
M31 218 216 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=102460 $D=1
M32 10 9 217 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=97830 $D=1
M33 11 9 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=102460 $D=1
M34 219 215 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=97830 $D=1
M35 220 216 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=102460 $D=1
M36 221 9 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=97830 $D=1
M37 222 9 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=102460 $D=1
M38 225 215 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=97830 $D=1
M39 226 216 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=102460 $D=1
M40 213 9 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=97830 $D=1
M41 214 9 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=102460 $D=1
M42 229 227 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=97830 $D=1
M43 230 228 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=102460 $D=1
M44 227 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=97830 $D=1
M45 228 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=102460 $D=1
M46 231 227 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=97830 $D=1
M47 232 228 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=102460 $D=1
M48 217 14 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=97830 $D=1
M49 218 14 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=102460 $D=1
M50 233 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=97830 $D=1
M51 234 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=102460 $D=1
M52 235 233 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=97830 $D=1
M53 236 234 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=102460 $D=1
M54 229 15 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=97830 $D=1
M55 230 15 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=102460 $D=1
M56 5 16 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=97830 $D=1
M57 6 16 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=102460 $D=1
M58 239 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=97830 $D=1
M59 240 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=102460 $D=1
M60 241 16 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=97830 $D=1
M61 242 16 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=102460 $D=1
M62 5 241 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=97830 $D=1
M63 6 242 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=102460 $D=1
M64 243 707 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=97830 $D=1
M65 244 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=102460 $D=1
M66 241 237 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=97830 $D=1
M67 242 238 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=102460 $D=1
M68 243 17 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=97830 $D=1
M69 244 17 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=102460 $D=1
M70 249 18 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=97830 $D=1
M71 250 18 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=102460 $D=1
M72 247 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=97830 $D=1
M73 248 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=102460 $D=1
M74 5 19 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=97830 $D=1
M75 6 19 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=102460 $D=1
M76 253 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=97830 $D=1
M77 254 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=102460 $D=1
M78 255 19 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=97830 $D=1
M79 256 19 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=102460 $D=1
M80 5 255 709 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=97830 $D=1
M81 6 256 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=102460 $D=1
M82 257 709 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=97830 $D=1
M83 258 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=102460 $D=1
M84 255 251 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=97830 $D=1
M85 256 252 258 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=102460 $D=1
M86 257 20 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=97830 $D=1
M87 258 20 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=102460 $D=1
M88 249 21 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=97830 $D=1
M89 250 21 258 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=102460 $D=1
M90 259 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=97830 $D=1
M91 260 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=102460 $D=1
M92 5 22 261 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=97830 $D=1
M93 6 22 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=102460 $D=1
M94 263 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=97830 $D=1
M95 264 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=102460 $D=1
M96 265 22 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=97830 $D=1
M97 266 22 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=102460 $D=1
M98 5 265 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=97830 $D=1
M99 6 266 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=102460 $D=1
M100 267 711 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=97830 $D=1
M101 268 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=102460 $D=1
M102 265 261 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=97830 $D=1
M103 266 262 268 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=102460 $D=1
M104 267 23 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=97830 $D=1
M105 268 23 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=102460 $D=1
M106 249 24 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=97830 $D=1
M107 250 24 268 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=102460 $D=1
M108 269 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=97830 $D=1
M109 270 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=102460 $D=1
M110 5 25 271 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=97830 $D=1
M111 6 25 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=102460 $D=1
M112 273 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=97830 $D=1
M113 274 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=102460 $D=1
M114 275 25 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=97830 $D=1
M115 276 25 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=102460 $D=1
M116 5 275 713 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=97830 $D=1
M117 6 276 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=102460 $D=1
M118 277 713 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=97830 $D=1
M119 278 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=102460 $D=1
M120 275 271 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=97830 $D=1
M121 276 272 278 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=102460 $D=1
M122 277 26 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=97830 $D=1
M123 278 26 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=102460 $D=1
M124 249 27 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=97830 $D=1
M125 250 27 278 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=102460 $D=1
M126 279 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=97830 $D=1
M127 280 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=102460 $D=1
M128 5 28 281 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=97830 $D=1
M129 6 28 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=102460 $D=1
M130 283 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=97830 $D=1
M131 284 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=102460 $D=1
M132 285 28 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=97830 $D=1
M133 286 28 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=102460 $D=1
M134 5 285 715 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=97830 $D=1
M135 6 286 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=102460 $D=1
M136 287 715 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=97830 $D=1
M137 288 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=102460 $D=1
M138 285 281 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=97830 $D=1
M139 286 282 288 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=102460 $D=1
M140 287 29 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=97830 $D=1
M141 288 29 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=102460 $D=1
M142 249 30 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=97830 $D=1
M143 250 30 288 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=102460 $D=1
M144 289 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=97830 $D=1
M145 290 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=102460 $D=1
M146 5 31 291 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=97830 $D=1
M147 6 31 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=102460 $D=1
M148 293 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=97830 $D=1
M149 294 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=102460 $D=1
M150 295 31 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=97830 $D=1
M151 296 31 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=102460 $D=1
M152 5 295 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=97830 $D=1
M153 6 296 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=102460 $D=1
M154 297 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=97830 $D=1
M155 298 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=102460 $D=1
M156 295 291 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=97830 $D=1
M157 296 292 298 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=102460 $D=1
M158 297 32 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=97830 $D=1
M159 298 32 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=102460 $D=1
M160 249 33 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=97830 $D=1
M161 250 33 298 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=102460 $D=1
M162 299 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=97830 $D=1
M163 300 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=102460 $D=1
M164 5 34 301 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=97830 $D=1
M165 6 34 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=102460 $D=1
M166 303 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=97830 $D=1
M167 304 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=102460 $D=1
M168 305 34 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=97830 $D=1
M169 306 34 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=102460 $D=1
M170 5 305 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=97830 $D=1
M171 6 306 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=102460 $D=1
M172 307 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=97830 $D=1
M173 308 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=102460 $D=1
M174 305 301 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=97830 $D=1
M175 306 302 308 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=102460 $D=1
M176 307 35 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=97830 $D=1
M177 308 35 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=102460 $D=1
M178 249 36 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=97830 $D=1
M179 250 36 308 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=102460 $D=1
M180 309 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=97830 $D=1
M181 310 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=102460 $D=1
M182 5 37 311 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=97830 $D=1
M183 6 37 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=102460 $D=1
M184 313 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=97830 $D=1
M185 314 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=102460 $D=1
M186 315 37 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=97830 $D=1
M187 316 37 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=102460 $D=1
M188 5 315 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=97830 $D=1
M189 6 316 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=102460 $D=1
M190 317 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=97830 $D=1
M191 318 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=102460 $D=1
M192 315 311 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=97830 $D=1
M193 316 312 318 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=102460 $D=1
M194 317 38 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=97830 $D=1
M195 318 38 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=102460 $D=1
M196 249 39 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=97830 $D=1
M197 250 39 318 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=102460 $D=1
M198 319 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=97830 $D=1
M199 320 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=102460 $D=1
M200 5 40 321 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=97830 $D=1
M201 6 40 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=102460 $D=1
M202 323 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=97830 $D=1
M203 324 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=102460 $D=1
M204 325 40 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=97830 $D=1
M205 326 40 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=102460 $D=1
M206 5 325 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=97830 $D=1
M207 6 326 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=102460 $D=1
M208 327 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=97830 $D=1
M209 328 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=102460 $D=1
M210 325 321 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=97830 $D=1
M211 326 322 328 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=102460 $D=1
M212 327 41 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=97830 $D=1
M213 328 41 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=102460 $D=1
M214 249 42 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=97830 $D=1
M215 250 42 328 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=102460 $D=1
M216 329 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=97830 $D=1
M217 330 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=102460 $D=1
M218 5 43 331 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=97830 $D=1
M219 6 43 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=102460 $D=1
M220 333 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=97830 $D=1
M221 334 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=102460 $D=1
M222 335 43 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=97830 $D=1
M223 336 43 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=102460 $D=1
M224 5 335 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=97830 $D=1
M225 6 336 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=102460 $D=1
M226 337 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=97830 $D=1
M227 338 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=102460 $D=1
M228 335 331 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=97830 $D=1
M229 336 332 338 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=102460 $D=1
M230 337 44 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=97830 $D=1
M231 338 44 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=102460 $D=1
M232 249 45 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=97830 $D=1
M233 250 45 338 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=102460 $D=1
M234 339 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=97830 $D=1
M235 340 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=102460 $D=1
M236 5 46 341 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=97830 $D=1
M237 6 46 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=102460 $D=1
M238 343 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=97830 $D=1
M239 344 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=102460 $D=1
M240 345 46 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=97830 $D=1
M241 346 46 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=102460 $D=1
M242 5 345 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=97830 $D=1
M243 6 346 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=102460 $D=1
M244 347 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=97830 $D=1
M245 348 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=102460 $D=1
M246 345 341 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=97830 $D=1
M247 346 342 348 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=102460 $D=1
M248 347 47 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=97830 $D=1
M249 348 47 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=102460 $D=1
M250 249 48 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=97830 $D=1
M251 250 48 348 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=102460 $D=1
M252 349 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=97830 $D=1
M253 350 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=102460 $D=1
M254 5 49 351 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=97830 $D=1
M255 6 49 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=102460 $D=1
M256 353 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=97830 $D=1
M257 354 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=102460 $D=1
M258 355 49 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=97830 $D=1
M259 356 49 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=102460 $D=1
M260 5 355 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=97830 $D=1
M261 6 356 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=102460 $D=1
M262 357 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=97830 $D=1
M263 358 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=102460 $D=1
M264 355 351 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=97830 $D=1
M265 356 352 358 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=102460 $D=1
M266 357 50 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=97830 $D=1
M267 358 50 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=102460 $D=1
M268 249 51 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=97830 $D=1
M269 250 51 358 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=102460 $D=1
M270 359 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=97830 $D=1
M271 360 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=102460 $D=1
M272 5 52 361 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=97830 $D=1
M273 6 52 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=102460 $D=1
M274 363 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=97830 $D=1
M275 364 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=102460 $D=1
M276 365 52 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=97830 $D=1
M277 366 52 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=102460 $D=1
M278 5 365 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=97830 $D=1
M279 6 366 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=102460 $D=1
M280 367 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=97830 $D=1
M281 368 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=102460 $D=1
M282 365 361 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=97830 $D=1
M283 366 362 368 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=102460 $D=1
M284 367 53 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=97830 $D=1
M285 368 53 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=102460 $D=1
M286 249 54 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=97830 $D=1
M287 250 54 368 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=102460 $D=1
M288 369 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=97830 $D=1
M289 370 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=102460 $D=1
M290 5 55 371 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=97830 $D=1
M291 6 55 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=102460 $D=1
M292 373 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=97830 $D=1
M293 374 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=102460 $D=1
M294 375 55 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=97830 $D=1
M295 376 55 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=102460 $D=1
M296 5 375 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=97830 $D=1
M297 6 376 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=102460 $D=1
M298 377 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=97830 $D=1
M299 378 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=102460 $D=1
M300 375 371 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=97830 $D=1
M301 376 372 378 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=102460 $D=1
M302 377 56 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=97830 $D=1
M303 378 56 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=102460 $D=1
M304 249 57 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=97830 $D=1
M305 250 57 378 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=102460 $D=1
M306 379 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=97830 $D=1
M307 380 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=102460 $D=1
M308 5 58 381 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=97830 $D=1
M309 6 58 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=102460 $D=1
M310 383 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=97830 $D=1
M311 384 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=102460 $D=1
M312 385 58 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=97830 $D=1
M313 386 58 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=102460 $D=1
M314 5 385 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=97830 $D=1
M315 6 386 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=102460 $D=1
M316 387 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=97830 $D=1
M317 388 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=102460 $D=1
M318 385 381 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=97830 $D=1
M319 386 382 388 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=102460 $D=1
M320 387 59 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=97830 $D=1
M321 388 59 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=102460 $D=1
M322 249 60 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=97830 $D=1
M323 250 60 388 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=102460 $D=1
M324 389 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=97830 $D=1
M325 390 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=102460 $D=1
M326 5 61 391 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=97830 $D=1
M327 6 61 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=102460 $D=1
M328 393 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=97830 $D=1
M329 394 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=102460 $D=1
M330 395 61 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=97830 $D=1
M331 396 61 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=102460 $D=1
M332 5 395 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=97830 $D=1
M333 6 396 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=102460 $D=1
M334 397 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=97830 $D=1
M335 398 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=102460 $D=1
M336 395 391 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=97830 $D=1
M337 396 392 398 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=102460 $D=1
M338 397 62 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=97830 $D=1
M339 398 62 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=102460 $D=1
M340 249 63 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=97830 $D=1
M341 250 63 398 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=102460 $D=1
M342 399 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=97830 $D=1
M343 400 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=102460 $D=1
M344 5 64 401 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=97830 $D=1
M345 6 64 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=102460 $D=1
M346 403 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=97830 $D=1
M347 404 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=102460 $D=1
M348 405 64 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=97830 $D=1
M349 406 64 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=102460 $D=1
M350 5 405 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=97830 $D=1
M351 6 406 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=102460 $D=1
M352 407 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=97830 $D=1
M353 408 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=102460 $D=1
M354 405 401 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=97830 $D=1
M355 406 402 408 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=102460 $D=1
M356 407 65 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=97830 $D=1
M357 408 65 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=102460 $D=1
M358 249 66 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=97830 $D=1
M359 250 66 408 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=102460 $D=1
M360 409 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=97830 $D=1
M361 410 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=102460 $D=1
M362 5 67 411 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=97830 $D=1
M363 6 67 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=102460 $D=1
M364 413 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=97830 $D=1
M365 414 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=102460 $D=1
M366 415 67 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=97830 $D=1
M367 416 67 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=102460 $D=1
M368 5 415 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=97830 $D=1
M369 6 416 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=102460 $D=1
M370 417 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=97830 $D=1
M371 418 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=102460 $D=1
M372 415 411 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=97830 $D=1
M373 416 412 418 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=102460 $D=1
M374 417 68 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=97830 $D=1
M375 418 68 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=102460 $D=1
M376 249 69 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=97830 $D=1
M377 250 69 418 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=102460 $D=1
M378 419 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=97830 $D=1
M379 420 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=102460 $D=1
M380 5 70 421 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=97830 $D=1
M381 6 70 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=102460 $D=1
M382 423 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=97830 $D=1
M383 424 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=102460 $D=1
M384 425 70 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=97830 $D=1
M385 426 70 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=102460 $D=1
M386 5 425 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=97830 $D=1
M387 6 426 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=102460 $D=1
M388 427 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=97830 $D=1
M389 428 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=102460 $D=1
M390 425 421 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=97830 $D=1
M391 426 422 428 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=102460 $D=1
M392 427 71 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=97830 $D=1
M393 428 71 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=102460 $D=1
M394 249 72 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=97830 $D=1
M395 250 72 428 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=102460 $D=1
M396 429 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=97830 $D=1
M397 430 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=102460 $D=1
M398 5 73 431 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=97830 $D=1
M399 6 73 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=102460 $D=1
M400 433 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=97830 $D=1
M401 434 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=102460 $D=1
M402 435 73 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=97830 $D=1
M403 436 73 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=102460 $D=1
M404 5 435 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=97830 $D=1
M405 6 436 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=102460 $D=1
M406 437 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=97830 $D=1
M407 438 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=102460 $D=1
M408 435 431 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=97830 $D=1
M409 436 432 438 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=102460 $D=1
M410 437 74 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=97830 $D=1
M411 438 74 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=102460 $D=1
M412 249 75 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=97830 $D=1
M413 250 75 438 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=102460 $D=1
M414 439 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=97830 $D=1
M415 440 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=102460 $D=1
M416 5 76 441 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=97830 $D=1
M417 6 76 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=102460 $D=1
M418 443 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=97830 $D=1
M419 444 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=102460 $D=1
M420 445 76 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=97830 $D=1
M421 446 76 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=102460 $D=1
M422 5 445 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=97830 $D=1
M423 6 446 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=102460 $D=1
M424 447 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=97830 $D=1
M425 448 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=102460 $D=1
M426 445 441 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=97830 $D=1
M427 446 442 448 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=102460 $D=1
M428 447 77 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=97830 $D=1
M429 448 77 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=102460 $D=1
M430 249 78 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=97830 $D=1
M431 250 78 448 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=102460 $D=1
M432 449 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=97830 $D=1
M433 450 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=102460 $D=1
M434 5 79 451 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=97830 $D=1
M435 6 79 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=102460 $D=1
M436 453 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=97830 $D=1
M437 454 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=102460 $D=1
M438 455 79 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=97830 $D=1
M439 456 79 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=102460 $D=1
M440 5 455 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=97830 $D=1
M441 6 456 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=102460 $D=1
M442 457 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=97830 $D=1
M443 458 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=102460 $D=1
M444 455 451 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=97830 $D=1
M445 456 452 458 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=102460 $D=1
M446 457 80 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=97830 $D=1
M447 458 80 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=102460 $D=1
M448 249 81 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=97830 $D=1
M449 250 81 458 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=102460 $D=1
M450 459 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=97830 $D=1
M451 460 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=102460 $D=1
M452 5 82 461 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=97830 $D=1
M453 6 82 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=102460 $D=1
M454 463 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=97830 $D=1
M455 464 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=102460 $D=1
M456 465 82 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=97830 $D=1
M457 466 82 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=102460 $D=1
M458 5 465 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=97830 $D=1
M459 6 466 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=102460 $D=1
M460 467 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=97830 $D=1
M461 468 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=102460 $D=1
M462 465 461 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=97830 $D=1
M463 466 462 468 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=102460 $D=1
M464 467 83 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=97830 $D=1
M465 468 83 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=102460 $D=1
M466 249 84 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=97830 $D=1
M467 250 84 468 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=102460 $D=1
M468 469 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=97830 $D=1
M469 470 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=102460 $D=1
M470 5 85 471 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=97830 $D=1
M471 6 85 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=102460 $D=1
M472 473 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=97830 $D=1
M473 474 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=102460 $D=1
M474 475 85 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=97830 $D=1
M475 476 85 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=102460 $D=1
M476 5 475 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=97830 $D=1
M477 6 476 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=102460 $D=1
M478 477 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=97830 $D=1
M479 478 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=102460 $D=1
M480 475 471 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=97830 $D=1
M481 476 472 478 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=102460 $D=1
M482 477 86 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=97830 $D=1
M483 478 86 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=102460 $D=1
M484 249 87 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=97830 $D=1
M485 250 87 478 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=102460 $D=1
M486 479 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=97830 $D=1
M487 480 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=102460 $D=1
M488 5 88 481 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=97830 $D=1
M489 6 88 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=102460 $D=1
M490 483 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=97830 $D=1
M491 484 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=102460 $D=1
M492 485 88 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=97830 $D=1
M493 486 88 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=102460 $D=1
M494 5 485 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=97830 $D=1
M495 6 486 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=102460 $D=1
M496 487 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=97830 $D=1
M497 488 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=102460 $D=1
M498 485 481 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=97830 $D=1
M499 486 482 488 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=102460 $D=1
M500 487 89 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=97830 $D=1
M501 488 89 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=102460 $D=1
M502 249 90 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=97830 $D=1
M503 250 90 488 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=102460 $D=1
M504 489 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=97830 $D=1
M505 490 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=102460 $D=1
M506 5 91 491 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=97830 $D=1
M507 6 91 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=102460 $D=1
M508 493 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=97830 $D=1
M509 494 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=102460 $D=1
M510 495 91 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=97830 $D=1
M511 496 91 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=102460 $D=1
M512 5 495 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=97830 $D=1
M513 6 496 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=102460 $D=1
M514 497 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=97830 $D=1
M515 498 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=102460 $D=1
M516 495 491 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=97830 $D=1
M517 496 492 498 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=102460 $D=1
M518 497 92 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=97830 $D=1
M519 498 92 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=102460 $D=1
M520 249 93 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=97830 $D=1
M521 250 93 498 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=102460 $D=1
M522 499 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=97830 $D=1
M523 500 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=102460 $D=1
M524 5 94 501 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=97830 $D=1
M525 6 94 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=102460 $D=1
M526 503 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=97830 $D=1
M527 504 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=102460 $D=1
M528 505 94 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=97830 $D=1
M529 506 94 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=102460 $D=1
M530 5 505 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=97830 $D=1
M531 6 506 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=102460 $D=1
M532 507 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=97830 $D=1
M533 508 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=102460 $D=1
M534 505 501 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=97830 $D=1
M535 506 502 508 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=102460 $D=1
M536 507 95 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=97830 $D=1
M537 508 95 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=102460 $D=1
M538 249 96 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=97830 $D=1
M539 250 96 508 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=102460 $D=1
M540 509 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=97830 $D=1
M541 510 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=102460 $D=1
M542 5 97 511 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=97830 $D=1
M543 6 97 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=102460 $D=1
M544 513 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=97830 $D=1
M545 514 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=102460 $D=1
M546 515 97 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=97830 $D=1
M547 516 97 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=102460 $D=1
M548 5 515 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=97830 $D=1
M549 6 516 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=102460 $D=1
M550 517 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=97830 $D=1
M551 518 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=102460 $D=1
M552 515 511 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=97830 $D=1
M553 516 512 518 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=102460 $D=1
M554 517 98 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=97830 $D=1
M555 518 98 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=102460 $D=1
M556 249 99 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=97830 $D=1
M557 250 99 518 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=102460 $D=1
M558 519 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=97830 $D=1
M559 520 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=102460 $D=1
M560 5 100 521 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=97830 $D=1
M561 6 100 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=102460 $D=1
M562 523 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=97830 $D=1
M563 524 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=102460 $D=1
M564 525 100 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=97830 $D=1
M565 526 100 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=102460 $D=1
M566 5 525 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=97830 $D=1
M567 6 526 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=102460 $D=1
M568 527 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=97830 $D=1
M569 528 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=102460 $D=1
M570 525 521 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=97830 $D=1
M571 526 522 528 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=102460 $D=1
M572 527 101 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=97830 $D=1
M573 528 101 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=102460 $D=1
M574 249 102 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=97830 $D=1
M575 250 102 528 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=102460 $D=1
M576 529 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=97830 $D=1
M577 530 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=102460 $D=1
M578 5 103 531 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=97830 $D=1
M579 6 103 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=102460 $D=1
M580 533 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=97830 $D=1
M581 534 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=102460 $D=1
M582 535 103 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=97830 $D=1
M583 536 103 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=102460 $D=1
M584 5 535 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=97830 $D=1
M585 6 536 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=102460 $D=1
M586 537 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=97830 $D=1
M587 538 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=102460 $D=1
M588 535 531 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=97830 $D=1
M589 536 532 538 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=102460 $D=1
M590 537 104 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=97830 $D=1
M591 538 104 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=102460 $D=1
M592 249 105 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=97830 $D=1
M593 250 105 538 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=102460 $D=1
M594 539 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=97830 $D=1
M595 540 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=102460 $D=1
M596 5 106 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=97830 $D=1
M597 6 106 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=102460 $D=1
M598 543 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=97830 $D=1
M599 544 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=102460 $D=1
M600 545 106 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=97830 $D=1
M601 546 106 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=102460 $D=1
M602 5 545 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=97830 $D=1
M603 6 546 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=102460 $D=1
M604 547 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=97830 $D=1
M605 548 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=102460 $D=1
M606 545 541 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=97830 $D=1
M607 546 542 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=102460 $D=1
M608 547 107 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=97830 $D=1
M609 548 107 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=102460 $D=1
M610 249 108 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=97830 $D=1
M611 250 108 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=102460 $D=1
M612 549 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=97830 $D=1
M613 550 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=102460 $D=1
M614 5 109 551 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=97830 $D=1
M615 6 109 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=102460 $D=1
M616 553 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=97830 $D=1
M617 554 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=102460 $D=1
M618 5 110 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=97830 $D=1
M619 6 110 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=102460 $D=1
M620 249 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=97830 $D=1
M621 250 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=102460 $D=1
M622 5 557 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=97830 $D=1
M623 6 558 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=102460 $D=1
M624 557 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=97830 $D=1
M625 558 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=102460 $D=1
M626 769 245 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=97830 $D=1
M627 770 246 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=102460 $D=1
M628 559 555 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=97830 $D=1
M629 560 556 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=102460 $D=1
M630 5 559 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=97830 $D=1
M631 6 560 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=102460 $D=1
M632 771 561 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=97830 $D=1
M633 772 562 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=102460 $D=1
M634 559 557 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=97830 $D=1
M635 560 558 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=102460 $D=1
M636 5 565 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=97830 $D=1
M637 6 566 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=102460 $D=1
M638 565 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=97830 $D=1
M639 566 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=102460 $D=1
M640 773 249 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=97830 $D=1
M641 774 250 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=102460 $D=1
M642 567 563 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=97830 $D=1
M643 568 564 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=102460 $D=1
M644 5 567 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=97830 $D=1
M645 6 568 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=102460 $D=1
M646 775 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=97830 $D=1
M647 776 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=102460 $D=1
M648 567 565 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=97830 $D=1
M649 568 566 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=102460 $D=1
M650 569 115 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=97830 $D=1
M651 570 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=102460 $D=1
M652 571 569 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=97830 $D=1
M653 572 570 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=102460 $D=1
M654 117 115 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=97830 $D=1
M655 117 115 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=102460 $D=1
M656 573 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=97830 $D=1
M657 574 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=102460 $D=1
M658 575 573 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=97830 $D=1
M659 576 574 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=102460 $D=1
M660 777 118 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=97830 $D=1
M661 778 118 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=102460 $D=1
M662 5 112 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=97830 $D=1
M663 6 113 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=102460 $D=1
M664 577 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=97830 $D=1
M665 578 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=102460 $D=1
M666 579 577 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=97830 $D=1
M667 580 578 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=102460 $D=1
M668 10 121 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=97830 $D=1
M669 11 121 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=102460 $D=1
M670 582 581 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=97830 $D=1
M671 583 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=102460 $D=1
M672 5 586 584 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=97830 $D=1
M673 6 587 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=102460 $D=1
M674 588 571 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=97830 $D=1
M675 589 572 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=102460 $D=1
M676 586 588 581 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=97830 $D=1
M677 587 589 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=102460 $D=1
M678 582 571 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=97830 $D=1
M679 583 572 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=102460 $D=1
M680 590 584 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=97830 $D=1
M681 591 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=102460 $D=1
M682 125 590 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=97830 $D=1
M683 581 591 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=102460 $D=1
M684 571 584 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=97830 $D=1
M685 572 585 581 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=102460 $D=1
M686 592 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=97830 $D=1
M687 593 581 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=102460 $D=1
M688 594 584 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=97830 $D=1
M689 595 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=102460 $D=1
M690 596 594 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=97830 $D=1
M691 597 595 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=102460 $D=1
M692 579 584 596 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=97830 $D=1
M693 580 585 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=102460 $D=1
M694 598 571 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=97830 $D=1
M695 599 572 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=102460 $D=1
M696 5 579 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=97830 $D=1
M697 6 580 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=102460 $D=1
M698 600 596 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=97830 $D=1
M699 601 597 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=102460 $D=1
M700 797 571 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=97830 $D=1
M701 798 572 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=102460 $D=1
M702 602 579 797 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=97830 $D=1
M703 603 580 798 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=102460 $D=1
M704 799 571 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=97830 $D=1
M705 800 572 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=102460 $D=1
M706 604 579 799 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=97830 $D=1
M707 605 580 800 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=102460 $D=1
M708 608 571 606 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=97830 $D=1
M709 609 572 607 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=102460 $D=1
M710 606 579 608 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=97830 $D=1
M711 607 580 609 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=102460 $D=1
M712 5 604 606 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=97830 $D=1
M713 6 605 607 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=102460 $D=1
M714 610 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=97830 $D=1
M715 611 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=102460 $D=1
M716 612 610 598 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=97830 $D=1
M717 613 611 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=102460 $D=1
M718 602 127 612 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=97830 $D=1
M719 603 127 613 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=102460 $D=1
M720 614 610 600 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=97830 $D=1
M721 615 611 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=102460 $D=1
M722 608 127 614 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=97830 $D=1
M723 609 127 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=102460 $D=1
M724 616 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=97830 $D=1
M725 617 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=102460 $D=1
M726 618 616 614 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=97830 $D=1
M727 619 617 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=102460 $D=1
M728 612 128 618 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=97830 $D=1
M729 613 128 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=102460 $D=1
M730 12 618 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=97830 $D=1
M731 13 619 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=102460 $D=1
M732 620 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=97830 $D=1
M733 621 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=102460 $D=1
M734 622 620 130 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=97830 $D=1
M735 623 621 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=102460 $D=1
M736 132 129 622 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=97830 $D=1
M737 133 129 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=102460 $D=1
M738 624 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=97830 $D=1
M739 625 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=102460 $D=1
M740 626 624 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=97830 $D=1
M741 627 625 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=102460 $D=1
M742 136 129 626 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=97830 $D=1
M743 137 129 627 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=102460 $D=1
M744 628 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=97830 $D=1
M745 629 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=102460 $D=1
M746 123 628 137 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=97830 $D=1
M747 123 629 138 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=102460 $D=1
M748 116 129 123 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=97830 $D=1
M749 120 129 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=102460 $D=1
M750 630 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=97830 $D=1
M751 631 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=102460 $D=1
M752 632 630 139 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=97830 $D=1
M753 633 631 140 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=102460 $D=1
M754 114 129 632 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=97830 $D=1
M755 119 129 633 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=102460 $D=1
M756 634 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=97830 $D=1
M757 635 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=102460 $D=1
M758 636 634 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=97830 $D=1
M759 637 635 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=102460 $D=1
M760 141 129 636 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=97830 $D=1
M761 142 129 637 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=102460 $D=1
M762 5 571 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=97830 $D=1
M763 6 572 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=102460 $D=1
M764 133 779 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=97830 $D=1
M765 130 780 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=102460 $D=1
M766 638 143 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=97830 $D=1
M767 639 143 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=102460 $D=1
M768 144 638 133 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=97830 $D=1
M769 145 639 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=102460 $D=1
M770 622 143 144 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=97830 $D=1
M771 623 143 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=102460 $D=1
M772 640 146 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=97830 $D=1
M773 641 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=102460 $D=1
M774 147 640 144 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=97830 $D=1
M775 126 641 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=102460 $D=1
M776 626 146 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=97830 $D=1
M777 627 146 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=102460 $D=1
M778 642 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=97830 $D=1
M779 643 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=102460 $D=1
M780 123 642 147 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=97830 $D=1
M781 124 643 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=102460 $D=1
M782 123 148 123 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=97830 $D=1
M783 123 148 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=102460 $D=1
M784 644 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=97830 $D=1
M785 645 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=102460 $D=1
M786 150 644 123 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=97830 $D=1
M787 151 645 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=102460 $D=1
M788 632 149 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=97830 $D=1
M789 633 149 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=102460 $D=1
M790 646 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=97830 $D=1
M791 647 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=102460 $D=1
M792 221 646 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=97830 $D=1
M793 222 647 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=102460 $D=1
M794 636 152 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=97830 $D=1
M795 637 152 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=102460 $D=1
M796 648 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=97830 $D=1
M797 649 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=102460 $D=1
M798 650 648 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=97830 $D=1
M799 651 649 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=102460 $D=1
M800 10 153 650 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=97830 $D=1
M801 11 153 651 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=102460 $D=1
M802 801 561 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=97830 $D=1
M803 802 562 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=102460 $D=1
M804 652 650 801 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=97830 $D=1
M805 653 651 802 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=102460 $D=1
M806 656 561 654 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=97830 $D=1
M807 657 562 655 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=102460 $D=1
M808 654 650 656 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=97830 $D=1
M809 655 651 657 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=102460 $D=1
M810 5 652 654 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=97830 $D=1
M811 6 653 655 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=102460 $D=1
M812 803 154 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=97830 $D=1
M813 804 658 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=102460 $D=1
M814 781 656 803 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=97830 $D=1
M815 782 657 804 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=102460 $D=1
M816 658 781 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=97830 $D=1
M817 155 782 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=102460 $D=1
M818 659 561 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=97830 $D=1
M819 660 562 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=102460 $D=1
M820 5 661 659 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=97830 $D=1
M821 6 662 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=102460 $D=1
M822 661 650 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=97830 $D=1
M823 662 651 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=102460 $D=1
M824 805 659 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=97830 $D=1
M825 806 660 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=102460 $D=1
M826 663 154 805 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=97830 $D=1
M827 664 658 806 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=102460 $D=1
M828 666 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=97830 $D=1
M829 667 665 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=102460 $D=1
M830 807 663 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=97830 $D=1
M831 808 664 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=102460 $D=1
M832 665 666 807 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=97830 $D=1
M833 157 667 808 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=102460 $D=1
M834 669 668 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=97830 $D=1
M835 670 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=102460 $D=1
M836 5 673 671 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=97830 $D=1
M837 6 674 672 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=102460 $D=1
M838 675 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=97830 $D=1
M839 676 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=102460 $D=1
M840 673 675 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=97830 $D=1
M841 674 676 158 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=102460 $D=1
M842 669 117 673 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=97830 $D=1
M843 670 117 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=102460 $D=1
M844 677 671 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=97830 $D=1
M845 678 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=102460 $D=1
M846 159 677 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=97830 $D=1
M847 668 678 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=102460 $D=1
M848 117 671 159 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=97830 $D=1
M849 117 672 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=102460 $D=1
M850 679 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=97830 $D=1
M851 680 668 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=102460 $D=1
M852 681 671 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=97830 $D=1
M853 682 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=102460 $D=1
M854 223 681 679 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=97830 $D=1
M855 224 682 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=102460 $D=1
M856 5 671 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=97830 $D=1
M857 6 672 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=102460 $D=1
M858 683 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=97830 $D=1
M859 684 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=102460 $D=1
M860 685 683 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=97830 $D=1
M861 686 684 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=102460 $D=1
M862 12 160 685 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=97830 $D=1
M863 13 160 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=102460 $D=1
M864 687 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=97830 $D=1
M865 688 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=102460 $D=1
M866 161 687 685 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=97830 $D=1
M867 161 688 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=102460 $D=1
M868 5 161 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=97830 $D=1
M869 6 161 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=102460 $D=1
M870 689 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=97830 $D=1
M871 690 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=102460 $D=1
M872 5 689 691 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=97830 $D=1
M873 6 690 692 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=102460 $D=1
M874 693 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=97830 $D=1
M875 694 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=102460 $D=1
M876 695 689 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=97830 $D=1
M877 696 690 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=102460 $D=1
M878 5 695 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=97830 $D=1
M879 6 696 784 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=102460 $D=1
M880 697 783 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=97830 $D=1
M881 698 784 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=102460 $D=1
M882 695 691 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=97830 $D=1
M883 696 692 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=102460 $D=1
M884 699 111 697 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=97830 $D=1
M885 700 111 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=102460 $D=1
M886 5 703 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=97830 $D=1
M887 6 704 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=102460 $D=1
M888 703 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=97830 $D=1
M889 704 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=102460 $D=1
M890 785 699 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=97830 $D=1
M891 786 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=102460 $D=1
M892 705 701 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=97830 $D=1
M893 706 702 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=102460 $D=1
M894 5 705 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=97830 $D=1
M895 6 706 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=102460 $D=1
M896 787 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=97830 $D=1
M897 788 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=102460 $D=1
M898 705 703 787 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=97830 $D=1
M899 706 704 788 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=102460 $D=1
M900 197 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=99080 $D=0
M901 198 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=103710 $D=0
M902 199 1 2 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=99080 $D=0
M903 200 1 3 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=103710 $D=0
M904 5 197 199 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=99080 $D=0
M905 6 198 200 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=103710 $D=0
M906 201 1 4 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=99080 $D=0
M907 202 1 4 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=103710 $D=0
M908 2 197 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=99080 $D=0
M909 3 198 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=103710 $D=0
M910 203 1 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=99080 $D=0
M911 204 1 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=103710 $D=0
M912 2 197 203 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=99080 $D=0
M913 3 198 204 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=103710 $D=0
M914 207 7 203 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=99080 $D=0
M915 208 7 204 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=103710 $D=0
M916 205 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=99080 $D=0
M917 206 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=103710 $D=0
M918 209 7 201 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=99080 $D=0
M919 210 7 202 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=103710 $D=0
M920 199 205 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=99080 $D=0
M921 200 206 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=103710 $D=0
M922 211 8 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=99080 $D=0
M923 212 8 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=103710 $D=0
M924 213 8 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=99080 $D=0
M925 214 8 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=103710 $D=0
M926 207 211 213 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=99080 $D=0
M927 208 212 214 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=103710 $D=0
M928 215 9 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=99080 $D=0
M929 216 9 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=103710 $D=0
M930 217 9 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=99080 $D=0
M931 218 9 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=103710 $D=0
M932 10 215 217 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=99080 $D=0
M933 11 216 218 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=103710 $D=0
M934 219 9 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=99080 $D=0
M935 220 9 13 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=103710 $D=0
M936 221 215 219 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=99080 $D=0
M937 222 216 220 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=103710 $D=0
M938 225 9 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=99080 $D=0
M939 226 9 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=103710 $D=0
M940 213 215 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=99080 $D=0
M941 214 216 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=103710 $D=0
M942 229 14 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=99080 $D=0
M943 230 14 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=103710 $D=0
M944 227 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=99080 $D=0
M945 228 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=103710 $D=0
M946 231 14 219 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=99080 $D=0
M947 232 14 220 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=103710 $D=0
M948 217 227 231 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=99080 $D=0
M949 218 228 232 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=103710 $D=0
M950 233 15 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=99080 $D=0
M951 234 15 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=103710 $D=0
M952 235 15 231 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=99080 $D=0
M953 236 15 232 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=103710 $D=0
M954 229 233 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=99080 $D=0
M955 230 234 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=103710 $D=0
M956 162 16 237 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=99080 $D=0
M957 163 16 238 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=103710 $D=0
M958 239 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=99080 $D=0
M959 240 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=103710 $D=0
M960 241 237 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=99080 $D=0
M961 242 238 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=103710 $D=0
M962 162 241 707 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=99080 $D=0
M963 163 242 708 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=103710 $D=0
M964 243 707 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=99080 $D=0
M965 244 708 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=103710 $D=0
M966 241 16 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=99080 $D=0
M967 242 16 244 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=103710 $D=0
M968 243 239 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=99080 $D=0
M969 244 240 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=103710 $D=0
M970 249 247 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=99080 $D=0
M971 250 248 244 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=103710 $D=0
M972 247 18 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=99080 $D=0
M973 248 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=103710 $D=0
M974 162 19 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=99080 $D=0
M975 163 19 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=103710 $D=0
M976 253 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=99080 $D=0
M977 254 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=103710 $D=0
M978 255 251 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=99080 $D=0
M979 256 252 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=103710 $D=0
M980 162 255 709 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=99080 $D=0
M981 163 256 710 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=103710 $D=0
M982 257 709 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=99080 $D=0
M983 258 710 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=103710 $D=0
M984 255 19 257 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=99080 $D=0
M985 256 19 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=103710 $D=0
M986 257 253 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=99080 $D=0
M987 258 254 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=103710 $D=0
M988 249 259 257 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=99080 $D=0
M989 250 260 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=103710 $D=0
M990 259 21 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=99080 $D=0
M991 260 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=103710 $D=0
M992 162 22 261 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=99080 $D=0
M993 163 22 262 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=103710 $D=0
M994 263 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=99080 $D=0
M995 264 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=103710 $D=0
M996 265 261 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=99080 $D=0
M997 266 262 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=103710 $D=0
M998 162 265 711 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=99080 $D=0
M999 163 266 712 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=103710 $D=0
M1000 267 711 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=99080 $D=0
M1001 268 712 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=103710 $D=0
M1002 265 22 267 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=99080 $D=0
M1003 266 22 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=103710 $D=0
M1004 267 263 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=99080 $D=0
M1005 268 264 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=103710 $D=0
M1006 249 269 267 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=99080 $D=0
M1007 250 270 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=103710 $D=0
M1008 269 24 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=99080 $D=0
M1009 270 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=103710 $D=0
M1010 162 25 271 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=99080 $D=0
M1011 163 25 272 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=103710 $D=0
M1012 273 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=99080 $D=0
M1013 274 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=103710 $D=0
M1014 275 271 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=99080 $D=0
M1015 276 272 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=103710 $D=0
M1016 162 275 713 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=99080 $D=0
M1017 163 276 714 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=103710 $D=0
M1018 277 713 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=99080 $D=0
M1019 278 714 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=103710 $D=0
M1020 275 25 277 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=99080 $D=0
M1021 276 25 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=103710 $D=0
M1022 277 273 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=99080 $D=0
M1023 278 274 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=103710 $D=0
M1024 249 279 277 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=99080 $D=0
M1025 250 280 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=103710 $D=0
M1026 279 27 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=99080 $D=0
M1027 280 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=103710 $D=0
M1028 162 28 281 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=99080 $D=0
M1029 163 28 282 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=103710 $D=0
M1030 283 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=99080 $D=0
M1031 284 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=103710 $D=0
M1032 285 281 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=99080 $D=0
M1033 286 282 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=103710 $D=0
M1034 162 285 715 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=99080 $D=0
M1035 163 286 716 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=103710 $D=0
M1036 287 715 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=99080 $D=0
M1037 288 716 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=103710 $D=0
M1038 285 28 287 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=99080 $D=0
M1039 286 28 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=103710 $D=0
M1040 287 283 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=99080 $D=0
M1041 288 284 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=103710 $D=0
M1042 249 289 287 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=99080 $D=0
M1043 250 290 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=103710 $D=0
M1044 289 30 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=99080 $D=0
M1045 290 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=103710 $D=0
M1046 162 31 291 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=99080 $D=0
M1047 163 31 292 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=103710 $D=0
M1048 293 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=99080 $D=0
M1049 294 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=103710 $D=0
M1050 295 291 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=99080 $D=0
M1051 296 292 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=103710 $D=0
M1052 162 295 717 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=99080 $D=0
M1053 163 296 718 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=103710 $D=0
M1054 297 717 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=99080 $D=0
M1055 298 718 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=103710 $D=0
M1056 295 31 297 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=99080 $D=0
M1057 296 31 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=103710 $D=0
M1058 297 293 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=99080 $D=0
M1059 298 294 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=103710 $D=0
M1060 249 299 297 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=99080 $D=0
M1061 250 300 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=103710 $D=0
M1062 299 33 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=99080 $D=0
M1063 300 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=103710 $D=0
M1064 162 34 301 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=99080 $D=0
M1065 163 34 302 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=103710 $D=0
M1066 303 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=99080 $D=0
M1067 304 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=103710 $D=0
M1068 305 301 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=99080 $D=0
M1069 306 302 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=103710 $D=0
M1070 162 305 719 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=99080 $D=0
M1071 163 306 720 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=103710 $D=0
M1072 307 719 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=99080 $D=0
M1073 308 720 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=103710 $D=0
M1074 305 34 307 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=99080 $D=0
M1075 306 34 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=103710 $D=0
M1076 307 303 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=99080 $D=0
M1077 308 304 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=103710 $D=0
M1078 249 309 307 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=99080 $D=0
M1079 250 310 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=103710 $D=0
M1080 309 36 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=99080 $D=0
M1081 310 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=103710 $D=0
M1082 162 37 311 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=99080 $D=0
M1083 163 37 312 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=103710 $D=0
M1084 313 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=99080 $D=0
M1085 314 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=103710 $D=0
M1086 315 311 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=99080 $D=0
M1087 316 312 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=103710 $D=0
M1088 162 315 721 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=99080 $D=0
M1089 163 316 722 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=103710 $D=0
M1090 317 721 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=99080 $D=0
M1091 318 722 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=103710 $D=0
M1092 315 37 317 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=99080 $D=0
M1093 316 37 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=103710 $D=0
M1094 317 313 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=99080 $D=0
M1095 318 314 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=103710 $D=0
M1096 249 319 317 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=99080 $D=0
M1097 250 320 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=103710 $D=0
M1098 319 39 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=99080 $D=0
M1099 320 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=103710 $D=0
M1100 162 40 321 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=99080 $D=0
M1101 163 40 322 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=103710 $D=0
M1102 323 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=99080 $D=0
M1103 324 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=103710 $D=0
M1104 325 321 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=99080 $D=0
M1105 326 322 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=103710 $D=0
M1106 162 325 723 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=99080 $D=0
M1107 163 326 724 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=103710 $D=0
M1108 327 723 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=99080 $D=0
M1109 328 724 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=103710 $D=0
M1110 325 40 327 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=99080 $D=0
M1111 326 40 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=103710 $D=0
M1112 327 323 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=99080 $D=0
M1113 328 324 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=103710 $D=0
M1114 249 329 327 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=99080 $D=0
M1115 250 330 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=103710 $D=0
M1116 329 42 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=99080 $D=0
M1117 330 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=103710 $D=0
M1118 162 43 331 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=99080 $D=0
M1119 163 43 332 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=103710 $D=0
M1120 333 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=99080 $D=0
M1121 334 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=103710 $D=0
M1122 335 331 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=99080 $D=0
M1123 336 332 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=103710 $D=0
M1124 162 335 725 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=99080 $D=0
M1125 163 336 726 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=103710 $D=0
M1126 337 725 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=99080 $D=0
M1127 338 726 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=103710 $D=0
M1128 335 43 337 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=99080 $D=0
M1129 336 43 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=103710 $D=0
M1130 337 333 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=99080 $D=0
M1131 338 334 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=103710 $D=0
M1132 249 339 337 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=99080 $D=0
M1133 250 340 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=103710 $D=0
M1134 339 45 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=99080 $D=0
M1135 340 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=103710 $D=0
M1136 162 46 341 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=99080 $D=0
M1137 163 46 342 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=103710 $D=0
M1138 343 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=99080 $D=0
M1139 344 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=103710 $D=0
M1140 345 341 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=99080 $D=0
M1141 346 342 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=103710 $D=0
M1142 162 345 727 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=99080 $D=0
M1143 163 346 728 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=103710 $D=0
M1144 347 727 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=99080 $D=0
M1145 348 728 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=103710 $D=0
M1146 345 46 347 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=99080 $D=0
M1147 346 46 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=103710 $D=0
M1148 347 343 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=99080 $D=0
M1149 348 344 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=103710 $D=0
M1150 249 349 347 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=99080 $D=0
M1151 250 350 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=103710 $D=0
M1152 349 48 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=99080 $D=0
M1153 350 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=103710 $D=0
M1154 162 49 351 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=99080 $D=0
M1155 163 49 352 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=103710 $D=0
M1156 353 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=99080 $D=0
M1157 354 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=103710 $D=0
M1158 355 351 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=99080 $D=0
M1159 356 352 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=103710 $D=0
M1160 162 355 729 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=99080 $D=0
M1161 163 356 730 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=103710 $D=0
M1162 357 729 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=99080 $D=0
M1163 358 730 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=103710 $D=0
M1164 355 49 357 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=99080 $D=0
M1165 356 49 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=103710 $D=0
M1166 357 353 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=99080 $D=0
M1167 358 354 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=103710 $D=0
M1168 249 359 357 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=99080 $D=0
M1169 250 360 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=103710 $D=0
M1170 359 51 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=99080 $D=0
M1171 360 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=103710 $D=0
M1172 162 52 361 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=99080 $D=0
M1173 163 52 362 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=103710 $D=0
M1174 363 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=99080 $D=0
M1175 364 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=103710 $D=0
M1176 365 361 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=99080 $D=0
M1177 366 362 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=103710 $D=0
M1178 162 365 731 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=99080 $D=0
M1179 163 366 732 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=103710 $D=0
M1180 367 731 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=99080 $D=0
M1181 368 732 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=103710 $D=0
M1182 365 52 367 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=99080 $D=0
M1183 366 52 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=103710 $D=0
M1184 367 363 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=99080 $D=0
M1185 368 364 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=103710 $D=0
M1186 249 369 367 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=99080 $D=0
M1187 250 370 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=103710 $D=0
M1188 369 54 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=99080 $D=0
M1189 370 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=103710 $D=0
M1190 162 55 371 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=99080 $D=0
M1191 163 55 372 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=103710 $D=0
M1192 373 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=99080 $D=0
M1193 374 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=103710 $D=0
M1194 375 371 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=99080 $D=0
M1195 376 372 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=103710 $D=0
M1196 162 375 733 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=99080 $D=0
M1197 163 376 734 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=103710 $D=0
M1198 377 733 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=99080 $D=0
M1199 378 734 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=103710 $D=0
M1200 375 55 377 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=99080 $D=0
M1201 376 55 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=103710 $D=0
M1202 377 373 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=99080 $D=0
M1203 378 374 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=103710 $D=0
M1204 249 379 377 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=99080 $D=0
M1205 250 380 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=103710 $D=0
M1206 379 57 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=99080 $D=0
M1207 380 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=103710 $D=0
M1208 162 58 381 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=99080 $D=0
M1209 163 58 382 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=103710 $D=0
M1210 383 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=99080 $D=0
M1211 384 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=103710 $D=0
M1212 385 381 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=99080 $D=0
M1213 386 382 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=103710 $D=0
M1214 162 385 735 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=99080 $D=0
M1215 163 386 736 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=103710 $D=0
M1216 387 735 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=99080 $D=0
M1217 388 736 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=103710 $D=0
M1218 385 58 387 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=99080 $D=0
M1219 386 58 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=103710 $D=0
M1220 387 383 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=99080 $D=0
M1221 388 384 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=103710 $D=0
M1222 249 389 387 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=99080 $D=0
M1223 250 390 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=103710 $D=0
M1224 389 60 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=99080 $D=0
M1225 390 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=103710 $D=0
M1226 162 61 391 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=99080 $D=0
M1227 163 61 392 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=103710 $D=0
M1228 393 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=99080 $D=0
M1229 394 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=103710 $D=0
M1230 395 391 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=99080 $D=0
M1231 396 392 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=103710 $D=0
M1232 162 395 737 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=99080 $D=0
M1233 163 396 738 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=103710 $D=0
M1234 397 737 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=99080 $D=0
M1235 398 738 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=103710 $D=0
M1236 395 61 397 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=99080 $D=0
M1237 396 61 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=103710 $D=0
M1238 397 393 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=99080 $D=0
M1239 398 394 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=103710 $D=0
M1240 249 399 397 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=99080 $D=0
M1241 250 400 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=103710 $D=0
M1242 399 63 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=99080 $D=0
M1243 400 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=103710 $D=0
M1244 162 64 401 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=99080 $D=0
M1245 163 64 402 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=103710 $D=0
M1246 403 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=99080 $D=0
M1247 404 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=103710 $D=0
M1248 405 401 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=99080 $D=0
M1249 406 402 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=103710 $D=0
M1250 162 405 739 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=99080 $D=0
M1251 163 406 740 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=103710 $D=0
M1252 407 739 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=99080 $D=0
M1253 408 740 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=103710 $D=0
M1254 405 64 407 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=99080 $D=0
M1255 406 64 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=103710 $D=0
M1256 407 403 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=99080 $D=0
M1257 408 404 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=103710 $D=0
M1258 249 409 407 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=99080 $D=0
M1259 250 410 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=103710 $D=0
M1260 409 66 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=99080 $D=0
M1261 410 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=103710 $D=0
M1262 162 67 411 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=99080 $D=0
M1263 163 67 412 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=103710 $D=0
M1264 413 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=99080 $D=0
M1265 414 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=103710 $D=0
M1266 415 411 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=99080 $D=0
M1267 416 412 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=103710 $D=0
M1268 162 415 741 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=99080 $D=0
M1269 163 416 742 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=103710 $D=0
M1270 417 741 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=99080 $D=0
M1271 418 742 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=103710 $D=0
M1272 415 67 417 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=99080 $D=0
M1273 416 67 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=103710 $D=0
M1274 417 413 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=99080 $D=0
M1275 418 414 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=103710 $D=0
M1276 249 419 417 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=99080 $D=0
M1277 250 420 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=103710 $D=0
M1278 419 69 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=99080 $D=0
M1279 420 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=103710 $D=0
M1280 162 70 421 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=99080 $D=0
M1281 163 70 422 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=103710 $D=0
M1282 423 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=99080 $D=0
M1283 424 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=103710 $D=0
M1284 425 421 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=99080 $D=0
M1285 426 422 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=103710 $D=0
M1286 162 425 743 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=99080 $D=0
M1287 163 426 744 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=103710 $D=0
M1288 427 743 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=99080 $D=0
M1289 428 744 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=103710 $D=0
M1290 425 70 427 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=99080 $D=0
M1291 426 70 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=103710 $D=0
M1292 427 423 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=99080 $D=0
M1293 428 424 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=103710 $D=0
M1294 249 429 427 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=99080 $D=0
M1295 250 430 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=103710 $D=0
M1296 429 72 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=99080 $D=0
M1297 430 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=103710 $D=0
M1298 162 73 431 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=99080 $D=0
M1299 163 73 432 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=103710 $D=0
M1300 433 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=99080 $D=0
M1301 434 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=103710 $D=0
M1302 435 431 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=99080 $D=0
M1303 436 432 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=103710 $D=0
M1304 162 435 745 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=99080 $D=0
M1305 163 436 746 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=103710 $D=0
M1306 437 745 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=99080 $D=0
M1307 438 746 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=103710 $D=0
M1308 435 73 437 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=99080 $D=0
M1309 436 73 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=103710 $D=0
M1310 437 433 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=99080 $D=0
M1311 438 434 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=103710 $D=0
M1312 249 439 437 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=99080 $D=0
M1313 250 440 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=103710 $D=0
M1314 439 75 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=99080 $D=0
M1315 440 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=103710 $D=0
M1316 162 76 441 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=99080 $D=0
M1317 163 76 442 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=103710 $D=0
M1318 443 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=99080 $D=0
M1319 444 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=103710 $D=0
M1320 445 441 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=99080 $D=0
M1321 446 442 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=103710 $D=0
M1322 162 445 747 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=99080 $D=0
M1323 163 446 748 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=103710 $D=0
M1324 447 747 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=99080 $D=0
M1325 448 748 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=103710 $D=0
M1326 445 76 447 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=99080 $D=0
M1327 446 76 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=103710 $D=0
M1328 447 443 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=99080 $D=0
M1329 448 444 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=103710 $D=0
M1330 249 449 447 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=99080 $D=0
M1331 250 450 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=103710 $D=0
M1332 449 78 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=99080 $D=0
M1333 450 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=103710 $D=0
M1334 162 79 451 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=99080 $D=0
M1335 163 79 452 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=103710 $D=0
M1336 453 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=99080 $D=0
M1337 454 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=103710 $D=0
M1338 455 451 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=99080 $D=0
M1339 456 452 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=103710 $D=0
M1340 162 455 749 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=99080 $D=0
M1341 163 456 750 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=103710 $D=0
M1342 457 749 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=99080 $D=0
M1343 458 750 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=103710 $D=0
M1344 455 79 457 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=99080 $D=0
M1345 456 79 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=103710 $D=0
M1346 457 453 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=99080 $D=0
M1347 458 454 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=103710 $D=0
M1348 249 459 457 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=99080 $D=0
M1349 250 460 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=103710 $D=0
M1350 459 81 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=99080 $D=0
M1351 460 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=103710 $D=0
M1352 162 82 461 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=99080 $D=0
M1353 163 82 462 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=103710 $D=0
M1354 463 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=99080 $D=0
M1355 464 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=103710 $D=0
M1356 465 461 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=99080 $D=0
M1357 466 462 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=103710 $D=0
M1358 162 465 751 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=99080 $D=0
M1359 163 466 752 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=103710 $D=0
M1360 467 751 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=99080 $D=0
M1361 468 752 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=103710 $D=0
M1362 465 82 467 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=99080 $D=0
M1363 466 82 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=103710 $D=0
M1364 467 463 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=99080 $D=0
M1365 468 464 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=103710 $D=0
M1366 249 469 467 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=99080 $D=0
M1367 250 470 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=103710 $D=0
M1368 469 84 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=99080 $D=0
M1369 470 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=103710 $D=0
M1370 162 85 471 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=99080 $D=0
M1371 163 85 472 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=103710 $D=0
M1372 473 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=99080 $D=0
M1373 474 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=103710 $D=0
M1374 475 471 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=99080 $D=0
M1375 476 472 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=103710 $D=0
M1376 162 475 753 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=99080 $D=0
M1377 163 476 754 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=103710 $D=0
M1378 477 753 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=99080 $D=0
M1379 478 754 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=103710 $D=0
M1380 475 85 477 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=99080 $D=0
M1381 476 85 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=103710 $D=0
M1382 477 473 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=99080 $D=0
M1383 478 474 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=103710 $D=0
M1384 249 479 477 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=99080 $D=0
M1385 250 480 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=103710 $D=0
M1386 479 87 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=99080 $D=0
M1387 480 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=103710 $D=0
M1388 162 88 481 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=99080 $D=0
M1389 163 88 482 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=103710 $D=0
M1390 483 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=99080 $D=0
M1391 484 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=103710 $D=0
M1392 485 481 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=99080 $D=0
M1393 486 482 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=103710 $D=0
M1394 162 485 755 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=99080 $D=0
M1395 163 486 756 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=103710 $D=0
M1396 487 755 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=99080 $D=0
M1397 488 756 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=103710 $D=0
M1398 485 88 487 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=99080 $D=0
M1399 486 88 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=103710 $D=0
M1400 487 483 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=99080 $D=0
M1401 488 484 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=103710 $D=0
M1402 249 489 487 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=99080 $D=0
M1403 250 490 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=103710 $D=0
M1404 489 90 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=99080 $D=0
M1405 490 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=103710 $D=0
M1406 162 91 491 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=99080 $D=0
M1407 163 91 492 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=103710 $D=0
M1408 493 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=99080 $D=0
M1409 494 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=103710 $D=0
M1410 495 491 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=99080 $D=0
M1411 496 492 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=103710 $D=0
M1412 162 495 757 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=99080 $D=0
M1413 163 496 758 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=103710 $D=0
M1414 497 757 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=99080 $D=0
M1415 498 758 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=103710 $D=0
M1416 495 91 497 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=99080 $D=0
M1417 496 91 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=103710 $D=0
M1418 497 493 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=99080 $D=0
M1419 498 494 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=103710 $D=0
M1420 249 499 497 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=99080 $D=0
M1421 250 500 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=103710 $D=0
M1422 499 93 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=99080 $D=0
M1423 500 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=103710 $D=0
M1424 162 94 501 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=99080 $D=0
M1425 163 94 502 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=103710 $D=0
M1426 503 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=99080 $D=0
M1427 504 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=103710 $D=0
M1428 505 501 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=99080 $D=0
M1429 506 502 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=103710 $D=0
M1430 162 505 759 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=99080 $D=0
M1431 163 506 760 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=103710 $D=0
M1432 507 759 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=99080 $D=0
M1433 508 760 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=103710 $D=0
M1434 505 94 507 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=99080 $D=0
M1435 506 94 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=103710 $D=0
M1436 507 503 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=99080 $D=0
M1437 508 504 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=103710 $D=0
M1438 249 509 507 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=99080 $D=0
M1439 250 510 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=103710 $D=0
M1440 509 96 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=99080 $D=0
M1441 510 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=103710 $D=0
M1442 162 97 511 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=99080 $D=0
M1443 163 97 512 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=103710 $D=0
M1444 513 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=99080 $D=0
M1445 514 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=103710 $D=0
M1446 515 511 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=99080 $D=0
M1447 516 512 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=103710 $D=0
M1448 162 515 761 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=99080 $D=0
M1449 163 516 762 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=103710 $D=0
M1450 517 761 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=99080 $D=0
M1451 518 762 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=103710 $D=0
M1452 515 97 517 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=99080 $D=0
M1453 516 97 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=103710 $D=0
M1454 517 513 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=99080 $D=0
M1455 518 514 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=103710 $D=0
M1456 249 519 517 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=99080 $D=0
M1457 250 520 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=103710 $D=0
M1458 519 99 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=99080 $D=0
M1459 520 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=103710 $D=0
M1460 162 100 521 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=99080 $D=0
M1461 163 100 522 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=103710 $D=0
M1462 523 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=99080 $D=0
M1463 524 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=103710 $D=0
M1464 525 521 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=99080 $D=0
M1465 526 522 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=103710 $D=0
M1466 162 525 763 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=99080 $D=0
M1467 163 526 764 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=103710 $D=0
M1468 527 763 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=99080 $D=0
M1469 528 764 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=103710 $D=0
M1470 525 100 527 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=99080 $D=0
M1471 526 100 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=103710 $D=0
M1472 527 523 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=99080 $D=0
M1473 528 524 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=103710 $D=0
M1474 249 529 527 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=99080 $D=0
M1475 250 530 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=103710 $D=0
M1476 529 102 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=99080 $D=0
M1477 530 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=103710 $D=0
M1478 162 103 531 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=99080 $D=0
M1479 163 103 532 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=103710 $D=0
M1480 533 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=99080 $D=0
M1481 534 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=103710 $D=0
M1482 535 531 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=99080 $D=0
M1483 536 532 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=103710 $D=0
M1484 162 535 765 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=99080 $D=0
M1485 163 536 766 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=103710 $D=0
M1486 537 765 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=99080 $D=0
M1487 538 766 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=103710 $D=0
M1488 535 103 537 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=99080 $D=0
M1489 536 103 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=103710 $D=0
M1490 537 533 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=99080 $D=0
M1491 538 534 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=103710 $D=0
M1492 249 539 537 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=99080 $D=0
M1493 250 540 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=103710 $D=0
M1494 539 105 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=99080 $D=0
M1495 540 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=103710 $D=0
M1496 162 106 541 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=99080 $D=0
M1497 163 106 542 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=103710 $D=0
M1498 543 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=99080 $D=0
M1499 544 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=103710 $D=0
M1500 545 541 235 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=99080 $D=0
M1501 546 542 236 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=103710 $D=0
M1502 162 545 767 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=99080 $D=0
M1503 163 546 768 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=103710 $D=0
M1504 547 767 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=99080 $D=0
M1505 548 768 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=103710 $D=0
M1506 545 106 547 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=99080 $D=0
M1507 546 106 548 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=103710 $D=0
M1508 547 543 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=99080 $D=0
M1509 548 544 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=103710 $D=0
M1510 249 549 547 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=99080 $D=0
M1511 250 550 548 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=103710 $D=0
M1512 549 108 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=99080 $D=0
M1513 550 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=103710 $D=0
M1514 162 109 551 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=99080 $D=0
M1515 163 109 552 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=103710 $D=0
M1516 553 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=99080 $D=0
M1517 554 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=103710 $D=0
M1518 5 553 245 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=99080 $D=0
M1519 6 554 246 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=103710 $D=0
M1520 249 551 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=99080 $D=0
M1521 250 552 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=103710 $D=0
M1522 162 557 555 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=99080 $D=0
M1523 163 558 556 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=103710 $D=0
M1524 557 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=99080 $D=0
M1525 558 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=103710 $D=0
M1526 769 245 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=99080 $D=0
M1527 770 246 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=103710 $D=0
M1528 559 557 769 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=99080 $D=0
M1529 560 558 770 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=103710 $D=0
M1530 162 559 561 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=99080 $D=0
M1531 163 560 562 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=103710 $D=0
M1532 771 561 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=99080 $D=0
M1533 772 562 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=103710 $D=0
M1534 559 555 771 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=99080 $D=0
M1535 560 556 772 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=103710 $D=0
M1536 162 565 563 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=99080 $D=0
M1537 163 566 564 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=103710 $D=0
M1538 565 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=99080 $D=0
M1539 566 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=103710 $D=0
M1540 773 249 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=99080 $D=0
M1541 774 250 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=103710 $D=0
M1542 567 565 773 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=99080 $D=0
M1543 568 566 774 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=103710 $D=0
M1544 162 567 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=99080 $D=0
M1545 163 568 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=103710 $D=0
M1546 775 112 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=99080 $D=0
M1547 776 113 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=103710 $D=0
M1548 567 563 775 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=99080 $D=0
M1549 568 564 776 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=103710 $D=0
M1550 569 115 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=99080 $D=0
M1551 570 115 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=103710 $D=0
M1552 571 115 561 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=99080 $D=0
M1553 572 115 562 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=103710 $D=0
M1554 117 569 571 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=99080 $D=0
M1555 117 570 572 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=103710 $D=0
M1556 573 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=99080 $D=0
M1557 574 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=103710 $D=0
M1558 575 118 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=99080 $D=0
M1559 576 118 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=103710 $D=0
M1560 777 573 575 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=99080 $D=0
M1561 778 574 576 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=103710 $D=0
M1562 162 112 777 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=99080 $D=0
M1563 163 113 778 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=103710 $D=0
M1564 577 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=99080 $D=0
M1565 578 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=103710 $D=0
M1566 579 121 575 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=99080 $D=0
M1567 580 121 576 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=103710 $D=0
M1568 10 577 579 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=99080 $D=0
M1569 11 578 580 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=103710 $D=0
M1570 582 581 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=99080 $D=0
M1571 583 122 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=103710 $D=0
M1572 162 586 584 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=99080 $D=0
M1573 163 587 585 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=103710 $D=0
M1574 588 571 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=99080 $D=0
M1575 589 572 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=103710 $D=0
M1576 586 571 581 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=99080 $D=0
M1577 587 572 122 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=103710 $D=0
M1578 582 588 586 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=99080 $D=0
M1579 583 589 587 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=103710 $D=0
M1580 590 584 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=99080 $D=0
M1581 591 585 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=103710 $D=0
M1582 125 584 579 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=99080 $D=0
M1583 581 585 580 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=103710 $D=0
M1584 571 590 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=99080 $D=0
M1585 572 591 581 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=103710 $D=0
M1586 592 125 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=99080 $D=0
M1587 593 581 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=103710 $D=0
M1588 594 584 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=99080 $D=0
M1589 595 585 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=103710 $D=0
M1590 596 584 592 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=99080 $D=0
M1591 597 585 593 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=103710 $D=0
M1592 579 594 596 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=99080 $D=0
M1593 580 595 597 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=103710 $D=0
M1594 789 571 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=98720 $D=0
M1595 790 572 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=103350 $D=0
M1596 598 579 789 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=98720 $D=0
M1597 599 580 790 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=103350 $D=0
M1598 600 596 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=99080 $D=0
M1599 601 597 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=103710 $D=0
M1600 602 571 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=99080 $D=0
M1601 603 572 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=103710 $D=0
M1602 162 579 602 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=99080 $D=0
M1603 163 580 603 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=103710 $D=0
M1604 604 571 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=99080 $D=0
M1605 605 572 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=103710 $D=0
M1606 162 579 604 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=99080 $D=0
M1607 163 580 605 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=103710 $D=0
M1608 791 571 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=98900 $D=0
M1609 792 572 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=103530 $D=0
M1610 608 579 791 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=98900 $D=0
M1611 609 580 792 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=103530 $D=0
M1612 162 604 608 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=99080 $D=0
M1613 163 605 609 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=103710 $D=0
M1614 610 127 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=99080 $D=0
M1615 611 127 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=103710 $D=0
M1616 612 127 598 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=99080 $D=0
M1617 613 127 599 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=103710 $D=0
M1618 602 610 612 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=99080 $D=0
M1619 603 611 613 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=103710 $D=0
M1620 614 127 600 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=99080 $D=0
M1621 615 127 601 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=103710 $D=0
M1622 608 610 614 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=99080 $D=0
M1623 609 611 615 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=103710 $D=0
M1624 616 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=99080 $D=0
M1625 617 128 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=103710 $D=0
M1626 618 128 614 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=99080 $D=0
M1627 619 128 615 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=103710 $D=0
M1628 612 616 618 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=99080 $D=0
M1629 613 617 619 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=103710 $D=0
M1630 12 618 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=99080 $D=0
M1631 13 619 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=103710 $D=0
M1632 620 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=99080 $D=0
M1633 621 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=103710 $D=0
M1634 622 129 130 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=99080 $D=0
M1635 623 129 131 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=103710 $D=0
M1636 132 620 622 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=99080 $D=0
M1637 133 621 623 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=103710 $D=0
M1638 624 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=99080 $D=0
M1639 625 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=103710 $D=0
M1640 626 129 134 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=99080 $D=0
M1641 627 129 135 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=103710 $D=0
M1642 136 624 626 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=99080 $D=0
M1643 137 625 627 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=103710 $D=0
M1644 628 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=99080 $D=0
M1645 629 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=103710 $D=0
M1646 123 129 137 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=99080 $D=0
M1647 123 129 138 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=103710 $D=0
M1648 116 628 123 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=99080 $D=0
M1649 120 629 123 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=103710 $D=0
M1650 630 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=99080 $D=0
M1651 631 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=103710 $D=0
M1652 632 129 139 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=99080 $D=0
M1653 633 129 140 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=103710 $D=0
M1654 114 630 632 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=99080 $D=0
M1655 119 631 633 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=103710 $D=0
M1656 634 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=99080 $D=0
M1657 635 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=103710 $D=0
M1658 636 129 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=99080 $D=0
M1659 637 129 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=103710 $D=0
M1660 141 634 636 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=99080 $D=0
M1661 142 635 637 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=103710 $D=0
M1662 162 571 779 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=99080 $D=0
M1663 163 572 780 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=103710 $D=0
M1664 133 779 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=99080 $D=0
M1665 130 780 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=103710 $D=0
M1666 638 143 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=99080 $D=0
M1667 639 143 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=103710 $D=0
M1668 144 143 133 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=99080 $D=0
M1669 145 143 130 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=103710 $D=0
M1670 622 638 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=99080 $D=0
M1671 623 639 145 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=103710 $D=0
M1672 640 146 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=99080 $D=0
M1673 641 146 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=103710 $D=0
M1674 147 146 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=99080 $D=0
M1675 126 146 145 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=103710 $D=0
M1676 626 640 147 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=99080 $D=0
M1677 627 641 126 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=103710 $D=0
M1678 642 148 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=99080 $D=0
M1679 643 148 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=103710 $D=0
M1680 123 148 147 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=99080 $D=0
M1681 124 148 126 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=103710 $D=0
M1682 123 642 123 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=99080 $D=0
M1683 123 643 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=103710 $D=0
M1684 644 149 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=99080 $D=0
M1685 645 149 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=103710 $D=0
M1686 150 149 123 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=99080 $D=0
M1687 151 149 124 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=103710 $D=0
M1688 632 644 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=99080 $D=0
M1689 633 645 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=103710 $D=0
M1690 646 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=99080 $D=0
M1691 647 152 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=103710 $D=0
M1692 221 152 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=99080 $D=0
M1693 222 152 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=103710 $D=0
M1694 636 646 221 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=99080 $D=0
M1695 637 647 222 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=103710 $D=0
M1696 648 153 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=99080 $D=0
M1697 649 153 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=103710 $D=0
M1698 650 153 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=99080 $D=0
M1699 651 153 113 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=103710 $D=0
M1700 10 648 650 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=99080 $D=0
M1701 11 649 651 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=103710 $D=0
M1702 652 561 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=99080 $D=0
M1703 653 562 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=103710 $D=0
M1704 162 650 652 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=99080 $D=0
M1705 163 651 653 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=103710 $D=0
M1706 793 561 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=98900 $D=0
M1707 794 562 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=103530 $D=0
M1708 656 650 793 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=98900 $D=0
M1709 657 651 794 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=103530 $D=0
M1710 162 652 656 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=99080 $D=0
M1711 163 653 657 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=103710 $D=0
M1712 781 154 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=99080 $D=0
M1713 782 658 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=103710 $D=0
M1714 162 656 781 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=99080 $D=0
M1715 163 657 782 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=103710 $D=0
M1716 658 781 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=99080 $D=0
M1717 155 782 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=103710 $D=0
M1718 795 561 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=98720 $D=0
M1719 796 562 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=103350 $D=0
M1720 659 661 795 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=98720 $D=0
M1721 660 662 796 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=103350 $D=0
M1722 661 650 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=99080 $D=0
M1723 662 651 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=103710 $D=0
M1724 663 659 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=99080 $D=0
M1725 664 660 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=103710 $D=0
M1726 162 154 663 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=99080 $D=0
M1727 163 658 664 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=103710 $D=0
M1728 666 156 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=99080 $D=0
M1729 667 665 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=103710 $D=0
M1730 665 663 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=99080 $D=0
M1731 157 664 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=103710 $D=0
M1732 162 666 665 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=99080 $D=0
M1733 163 667 157 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=103710 $D=0
M1734 669 668 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=99080 $D=0
M1735 670 158 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=103710 $D=0
M1736 162 673 671 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=99080 $D=0
M1737 163 674 672 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=103710 $D=0
M1738 675 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=99080 $D=0
M1739 676 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=103710 $D=0
M1740 673 117 668 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=99080 $D=0
M1741 674 117 158 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=103710 $D=0
M1742 669 675 673 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=99080 $D=0
M1743 670 676 674 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=103710 $D=0
M1744 677 671 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=99080 $D=0
M1745 678 672 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=103710 $D=0
M1746 159 671 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=99080 $D=0
M1747 668 672 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=103710 $D=0
M1748 117 677 159 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=99080 $D=0
M1749 117 678 668 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=103710 $D=0
M1750 679 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=99080 $D=0
M1751 680 668 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=103710 $D=0
M1752 681 671 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=99080 $D=0
M1753 682 672 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=103710 $D=0
M1754 223 671 679 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=99080 $D=0
M1755 224 672 680 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=103710 $D=0
M1756 5 681 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=99080 $D=0
M1757 6 682 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=103710 $D=0
M1758 683 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=99080 $D=0
M1759 684 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=103710 $D=0
M1760 685 160 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=99080 $D=0
M1761 686 160 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=103710 $D=0
M1762 12 683 685 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=99080 $D=0
M1763 13 684 686 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=103710 $D=0
M1764 687 161 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=99080 $D=0
M1765 688 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=103710 $D=0
M1766 161 161 685 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=99080 $D=0
M1767 161 161 686 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=103710 $D=0
M1768 5 687 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=99080 $D=0
M1769 6 688 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=103710 $D=0
M1770 689 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=99080 $D=0
M1771 690 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=103710 $D=0
M1772 162 689 691 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=99080 $D=0
M1773 163 690 692 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=103710 $D=0
M1774 693 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=99080 $D=0
M1775 694 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=103710 $D=0
M1776 695 691 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=99080 $D=0
M1777 696 692 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=103710 $D=0
M1778 162 695 783 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=99080 $D=0
M1779 163 696 784 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=103710 $D=0
M1780 697 783 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=99080 $D=0
M1781 698 784 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=103710 $D=0
M1782 695 689 697 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=99080 $D=0
M1783 696 690 698 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=103710 $D=0
M1784 699 693 697 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=99080 $D=0
M1785 700 694 698 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=103710 $D=0
M1786 162 703 701 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=99080 $D=0
M1787 163 704 702 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=103710 $D=0
M1788 703 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=99080 $D=0
M1789 704 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=103710 $D=0
M1790 785 699 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=99080 $D=0
M1791 786 700 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=103710 $D=0
M1792 705 703 785 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=99080 $D=0
M1793 706 704 786 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=103710 $D=0
M1794 162 705 117 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=99080 $D=0
M1795 163 706 117 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=103710 $D=0
M1796 787 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=99080 $D=0
M1797 788 117 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=103710 $D=0
M1798 705 701 787 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=99080 $D=0
M1799 706 702 788 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=103710 $D=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162
** N=815 EP=162 IP=1514 FDC=1800
M0 201 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=88570 $D=1
M1 202 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=93200 $D=1
M2 203 201 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=88570 $D=1
M3 204 202 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=93200 $D=1
M4 5 1 203 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=88570 $D=1
M5 6 1 204 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=93200 $D=1
M6 205 201 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=88570 $D=1
M7 206 202 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=93200 $D=1
M8 2 1 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=88570 $D=1
M9 3 1 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=93200 $D=1
M10 207 201 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=88570 $D=1
M11 208 202 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=93200 $D=1
M12 2 1 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=88570 $D=1
M13 3 1 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=93200 $D=1
M14 211 209 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=88570 $D=1
M15 212 210 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=93200 $D=1
M16 209 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=88570 $D=1
M17 210 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=93200 $D=1
M18 213 209 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=88570 $D=1
M19 214 210 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=93200 $D=1
M20 203 7 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=88570 $D=1
M21 204 7 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=93200 $D=1
M22 215 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=88570 $D=1
M23 216 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=93200 $D=1
M24 217 215 213 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=88570 $D=1
M25 218 216 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=93200 $D=1
M26 211 8 217 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=88570 $D=1
M27 212 8 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=93200 $D=1
M28 219 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=88570 $D=1
M29 220 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=93200 $D=1
M30 221 219 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=88570 $D=1
M31 222 220 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=93200 $D=1
M32 10 9 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=88570 $D=1
M33 11 9 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=93200 $D=1
M34 223 219 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=88570 $D=1
M35 224 220 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=93200 $D=1
M36 225 9 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=88570 $D=1
M37 226 9 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=93200 $D=1
M38 229 219 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=88570 $D=1
M39 230 220 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=93200 $D=1
M40 217 9 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=88570 $D=1
M41 218 9 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=93200 $D=1
M42 233 231 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=88570 $D=1
M43 234 232 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=93200 $D=1
M44 231 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=88570 $D=1
M45 232 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=93200 $D=1
M46 235 231 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=88570 $D=1
M47 236 232 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=93200 $D=1
M48 221 14 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=88570 $D=1
M49 222 14 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=93200 $D=1
M50 237 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=88570 $D=1
M51 238 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=93200 $D=1
M52 239 237 235 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=88570 $D=1
M53 240 238 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=93200 $D=1
M54 233 15 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=88570 $D=1
M55 234 15 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=93200 $D=1
M56 5 16 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=88570 $D=1
M57 6 16 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=93200 $D=1
M58 243 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=88570 $D=1
M59 244 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=93200 $D=1
M60 245 16 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=88570 $D=1
M61 246 16 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=93200 $D=1
M62 5 245 714 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=88570 $D=1
M63 6 246 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=93200 $D=1
M64 247 714 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=88570 $D=1
M65 248 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=93200 $D=1
M66 245 241 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=88570 $D=1
M67 246 242 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=93200 $D=1
M68 247 17 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=88570 $D=1
M69 248 17 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=93200 $D=1
M70 253 18 247 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=88570 $D=1
M71 254 18 248 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=93200 $D=1
M72 251 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=88570 $D=1
M73 252 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=93200 $D=1
M74 5 19 255 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=88570 $D=1
M75 6 19 256 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=93200 $D=1
M76 257 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=88570 $D=1
M77 258 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=93200 $D=1
M78 259 19 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=88570 $D=1
M79 260 19 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=93200 $D=1
M80 5 259 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=88570 $D=1
M81 6 260 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=93200 $D=1
M82 261 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=88570 $D=1
M83 262 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=93200 $D=1
M84 259 255 261 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=88570 $D=1
M85 260 256 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=93200 $D=1
M86 261 20 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=88570 $D=1
M87 262 20 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=93200 $D=1
M88 253 21 261 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=88570 $D=1
M89 254 21 262 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=93200 $D=1
M90 263 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=88570 $D=1
M91 264 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=93200 $D=1
M92 5 22 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=88570 $D=1
M93 6 22 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=93200 $D=1
M94 267 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=88570 $D=1
M95 268 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=93200 $D=1
M96 269 22 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=88570 $D=1
M97 270 22 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=93200 $D=1
M98 5 269 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=88570 $D=1
M99 6 270 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=93200 $D=1
M100 271 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=88570 $D=1
M101 272 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=93200 $D=1
M102 269 265 271 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=88570 $D=1
M103 270 266 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=93200 $D=1
M104 271 23 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=88570 $D=1
M105 272 23 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=93200 $D=1
M106 253 24 271 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=88570 $D=1
M107 254 24 272 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=93200 $D=1
M108 273 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=88570 $D=1
M109 274 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=93200 $D=1
M110 5 25 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=88570 $D=1
M111 6 25 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=93200 $D=1
M112 277 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=88570 $D=1
M113 278 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=93200 $D=1
M114 279 25 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=88570 $D=1
M115 280 25 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=93200 $D=1
M116 5 279 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=88570 $D=1
M117 6 280 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=93200 $D=1
M118 281 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=88570 $D=1
M119 282 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=93200 $D=1
M120 279 275 281 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=88570 $D=1
M121 280 276 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=93200 $D=1
M122 281 26 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=88570 $D=1
M123 282 26 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=93200 $D=1
M124 253 27 281 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=88570 $D=1
M125 254 27 282 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=93200 $D=1
M126 283 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=88570 $D=1
M127 284 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=93200 $D=1
M128 5 28 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=88570 $D=1
M129 6 28 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=93200 $D=1
M130 287 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=88570 $D=1
M131 288 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=93200 $D=1
M132 289 28 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=88570 $D=1
M133 290 28 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=93200 $D=1
M134 5 289 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=88570 $D=1
M135 6 290 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=93200 $D=1
M136 291 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=88570 $D=1
M137 292 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=93200 $D=1
M138 289 285 291 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=88570 $D=1
M139 290 286 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=93200 $D=1
M140 291 29 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=88570 $D=1
M141 292 29 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=93200 $D=1
M142 253 30 291 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=88570 $D=1
M143 254 30 292 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=93200 $D=1
M144 293 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=88570 $D=1
M145 294 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=93200 $D=1
M146 5 31 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=88570 $D=1
M147 6 31 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=93200 $D=1
M148 297 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=88570 $D=1
M149 298 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=93200 $D=1
M150 299 31 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=88570 $D=1
M151 300 31 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=93200 $D=1
M152 5 299 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=88570 $D=1
M153 6 300 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=93200 $D=1
M154 301 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=88570 $D=1
M155 302 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=93200 $D=1
M156 299 295 301 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=88570 $D=1
M157 300 296 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=93200 $D=1
M158 301 32 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=88570 $D=1
M159 302 32 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=93200 $D=1
M160 253 33 301 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=88570 $D=1
M161 254 33 302 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=93200 $D=1
M162 303 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=88570 $D=1
M163 304 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=93200 $D=1
M164 5 34 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=88570 $D=1
M165 6 34 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=93200 $D=1
M166 307 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=88570 $D=1
M167 308 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=93200 $D=1
M168 309 34 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=88570 $D=1
M169 310 34 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=93200 $D=1
M170 5 309 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=88570 $D=1
M171 6 310 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=93200 $D=1
M172 311 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=88570 $D=1
M173 312 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=93200 $D=1
M174 309 305 311 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=88570 $D=1
M175 310 306 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=93200 $D=1
M176 311 35 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=88570 $D=1
M177 312 35 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=93200 $D=1
M178 253 36 311 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=88570 $D=1
M179 254 36 312 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=93200 $D=1
M180 313 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=88570 $D=1
M181 314 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=93200 $D=1
M182 5 37 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=88570 $D=1
M183 6 37 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=93200 $D=1
M184 317 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=88570 $D=1
M185 318 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=93200 $D=1
M186 319 37 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=88570 $D=1
M187 320 37 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=93200 $D=1
M188 5 319 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=88570 $D=1
M189 6 320 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=93200 $D=1
M190 321 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=88570 $D=1
M191 322 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=93200 $D=1
M192 319 315 321 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=88570 $D=1
M193 320 316 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=93200 $D=1
M194 321 38 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=88570 $D=1
M195 322 38 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=93200 $D=1
M196 253 39 321 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=88570 $D=1
M197 254 39 322 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=93200 $D=1
M198 323 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=88570 $D=1
M199 324 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=93200 $D=1
M200 5 40 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=88570 $D=1
M201 6 40 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=93200 $D=1
M202 327 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=88570 $D=1
M203 328 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=93200 $D=1
M204 329 40 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=88570 $D=1
M205 330 40 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=93200 $D=1
M206 5 329 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=88570 $D=1
M207 6 330 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=93200 $D=1
M208 331 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=88570 $D=1
M209 332 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=93200 $D=1
M210 329 325 331 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=88570 $D=1
M211 330 326 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=93200 $D=1
M212 331 41 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=88570 $D=1
M213 332 41 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=93200 $D=1
M214 253 42 331 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=88570 $D=1
M215 254 42 332 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=93200 $D=1
M216 333 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=88570 $D=1
M217 334 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=93200 $D=1
M218 5 43 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=88570 $D=1
M219 6 43 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=93200 $D=1
M220 337 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=88570 $D=1
M221 338 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=93200 $D=1
M222 339 43 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=88570 $D=1
M223 340 43 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=93200 $D=1
M224 5 339 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=88570 $D=1
M225 6 340 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=93200 $D=1
M226 341 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=88570 $D=1
M227 342 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=93200 $D=1
M228 339 335 341 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=88570 $D=1
M229 340 336 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=93200 $D=1
M230 341 44 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=88570 $D=1
M231 342 44 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=93200 $D=1
M232 253 45 341 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=88570 $D=1
M233 254 45 342 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=93200 $D=1
M234 343 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=88570 $D=1
M235 344 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=93200 $D=1
M236 5 46 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=88570 $D=1
M237 6 46 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=93200 $D=1
M238 347 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=88570 $D=1
M239 348 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=93200 $D=1
M240 349 46 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=88570 $D=1
M241 350 46 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=93200 $D=1
M242 5 349 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=88570 $D=1
M243 6 350 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=93200 $D=1
M244 351 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=88570 $D=1
M245 352 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=93200 $D=1
M246 349 345 351 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=88570 $D=1
M247 350 346 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=93200 $D=1
M248 351 47 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=88570 $D=1
M249 352 47 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=93200 $D=1
M250 253 48 351 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=88570 $D=1
M251 254 48 352 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=93200 $D=1
M252 353 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=88570 $D=1
M253 354 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=93200 $D=1
M254 5 49 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=88570 $D=1
M255 6 49 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=93200 $D=1
M256 357 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=88570 $D=1
M257 358 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=93200 $D=1
M258 359 49 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=88570 $D=1
M259 360 49 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=93200 $D=1
M260 5 359 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=88570 $D=1
M261 6 360 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=93200 $D=1
M262 361 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=88570 $D=1
M263 362 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=93200 $D=1
M264 359 355 361 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=88570 $D=1
M265 360 356 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=93200 $D=1
M266 361 50 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=88570 $D=1
M267 362 50 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=93200 $D=1
M268 253 51 361 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=88570 $D=1
M269 254 51 362 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=93200 $D=1
M270 363 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=88570 $D=1
M271 364 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=93200 $D=1
M272 5 52 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=88570 $D=1
M273 6 52 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=93200 $D=1
M274 367 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=88570 $D=1
M275 368 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=93200 $D=1
M276 369 52 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=88570 $D=1
M277 370 52 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=93200 $D=1
M278 5 369 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=88570 $D=1
M279 6 370 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=93200 $D=1
M280 371 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=88570 $D=1
M281 372 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=93200 $D=1
M282 369 365 371 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=88570 $D=1
M283 370 366 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=93200 $D=1
M284 371 53 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=88570 $D=1
M285 372 53 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=93200 $D=1
M286 253 54 371 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=88570 $D=1
M287 254 54 372 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=93200 $D=1
M288 373 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=88570 $D=1
M289 374 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=93200 $D=1
M290 5 55 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=88570 $D=1
M291 6 55 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=93200 $D=1
M292 377 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=88570 $D=1
M293 378 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=93200 $D=1
M294 379 55 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=88570 $D=1
M295 380 55 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=93200 $D=1
M296 5 379 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=88570 $D=1
M297 6 380 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=93200 $D=1
M298 381 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=88570 $D=1
M299 382 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=93200 $D=1
M300 379 375 381 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=88570 $D=1
M301 380 376 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=93200 $D=1
M302 381 56 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=88570 $D=1
M303 382 56 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=93200 $D=1
M304 253 57 381 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=88570 $D=1
M305 254 57 382 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=93200 $D=1
M306 383 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=88570 $D=1
M307 384 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=93200 $D=1
M308 5 58 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=88570 $D=1
M309 6 58 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=93200 $D=1
M310 387 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=88570 $D=1
M311 388 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=93200 $D=1
M312 389 58 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=88570 $D=1
M313 390 58 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=93200 $D=1
M314 5 389 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=88570 $D=1
M315 6 390 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=93200 $D=1
M316 391 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=88570 $D=1
M317 392 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=93200 $D=1
M318 389 385 391 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=88570 $D=1
M319 390 386 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=93200 $D=1
M320 391 59 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=88570 $D=1
M321 392 59 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=93200 $D=1
M322 253 60 391 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=88570 $D=1
M323 254 60 392 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=93200 $D=1
M324 393 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=88570 $D=1
M325 394 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=93200 $D=1
M326 5 61 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=88570 $D=1
M327 6 61 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=93200 $D=1
M328 397 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=88570 $D=1
M329 398 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=93200 $D=1
M330 399 61 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=88570 $D=1
M331 400 61 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=93200 $D=1
M332 5 399 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=88570 $D=1
M333 6 400 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=93200 $D=1
M334 401 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=88570 $D=1
M335 402 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=93200 $D=1
M336 399 395 401 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=88570 $D=1
M337 400 396 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=93200 $D=1
M338 401 62 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=88570 $D=1
M339 402 62 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=93200 $D=1
M340 253 63 401 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=88570 $D=1
M341 254 63 402 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=93200 $D=1
M342 403 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=88570 $D=1
M343 404 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=93200 $D=1
M344 5 64 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=88570 $D=1
M345 6 64 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=93200 $D=1
M346 407 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=88570 $D=1
M347 408 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=93200 $D=1
M348 409 64 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=88570 $D=1
M349 410 64 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=93200 $D=1
M350 5 409 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=88570 $D=1
M351 6 410 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=93200 $D=1
M352 411 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=88570 $D=1
M353 412 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=93200 $D=1
M354 409 405 411 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=88570 $D=1
M355 410 406 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=93200 $D=1
M356 411 65 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=88570 $D=1
M357 412 65 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=93200 $D=1
M358 253 66 411 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=88570 $D=1
M359 254 66 412 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=93200 $D=1
M360 413 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=88570 $D=1
M361 414 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=93200 $D=1
M362 5 67 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=88570 $D=1
M363 6 67 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=93200 $D=1
M364 417 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=88570 $D=1
M365 418 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=93200 $D=1
M366 419 67 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=88570 $D=1
M367 420 67 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=93200 $D=1
M368 5 419 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=88570 $D=1
M369 6 420 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=93200 $D=1
M370 421 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=88570 $D=1
M371 422 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=93200 $D=1
M372 419 415 421 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=88570 $D=1
M373 420 416 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=93200 $D=1
M374 421 68 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=88570 $D=1
M375 422 68 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=93200 $D=1
M376 253 69 421 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=88570 $D=1
M377 254 69 422 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=93200 $D=1
M378 423 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=88570 $D=1
M379 424 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=93200 $D=1
M380 5 70 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=88570 $D=1
M381 6 70 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=93200 $D=1
M382 427 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=88570 $D=1
M383 428 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=93200 $D=1
M384 429 70 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=88570 $D=1
M385 430 70 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=93200 $D=1
M386 5 429 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=88570 $D=1
M387 6 430 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=93200 $D=1
M388 431 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=88570 $D=1
M389 432 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=93200 $D=1
M390 429 425 431 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=88570 $D=1
M391 430 426 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=93200 $D=1
M392 431 71 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=88570 $D=1
M393 432 71 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=93200 $D=1
M394 253 72 431 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=88570 $D=1
M395 254 72 432 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=93200 $D=1
M396 433 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=88570 $D=1
M397 434 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=93200 $D=1
M398 5 73 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=88570 $D=1
M399 6 73 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=93200 $D=1
M400 437 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=88570 $D=1
M401 438 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=93200 $D=1
M402 439 73 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=88570 $D=1
M403 440 73 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=93200 $D=1
M404 5 439 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=88570 $D=1
M405 6 440 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=93200 $D=1
M406 441 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=88570 $D=1
M407 442 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=93200 $D=1
M408 439 435 441 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=88570 $D=1
M409 440 436 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=93200 $D=1
M410 441 74 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=88570 $D=1
M411 442 74 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=93200 $D=1
M412 253 75 441 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=88570 $D=1
M413 254 75 442 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=93200 $D=1
M414 443 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=88570 $D=1
M415 444 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=93200 $D=1
M416 5 76 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=88570 $D=1
M417 6 76 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=93200 $D=1
M418 447 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=88570 $D=1
M419 448 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=93200 $D=1
M420 449 76 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=88570 $D=1
M421 450 76 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=93200 $D=1
M422 5 449 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=88570 $D=1
M423 6 450 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=93200 $D=1
M424 451 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=88570 $D=1
M425 452 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=93200 $D=1
M426 449 445 451 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=88570 $D=1
M427 450 446 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=93200 $D=1
M428 451 77 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=88570 $D=1
M429 452 77 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=93200 $D=1
M430 253 78 451 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=88570 $D=1
M431 254 78 452 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=93200 $D=1
M432 453 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=88570 $D=1
M433 454 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=93200 $D=1
M434 5 79 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=88570 $D=1
M435 6 79 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=93200 $D=1
M436 457 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=88570 $D=1
M437 458 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=93200 $D=1
M438 459 79 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=88570 $D=1
M439 460 79 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=93200 $D=1
M440 5 459 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=88570 $D=1
M441 6 460 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=93200 $D=1
M442 461 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=88570 $D=1
M443 462 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=93200 $D=1
M444 459 455 461 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=88570 $D=1
M445 460 456 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=93200 $D=1
M446 461 80 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=88570 $D=1
M447 462 80 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=93200 $D=1
M448 253 81 461 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=88570 $D=1
M449 254 81 462 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=93200 $D=1
M450 463 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=88570 $D=1
M451 464 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=93200 $D=1
M452 5 82 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=88570 $D=1
M453 6 82 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=93200 $D=1
M454 467 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=88570 $D=1
M455 468 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=93200 $D=1
M456 469 82 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=88570 $D=1
M457 470 82 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=93200 $D=1
M458 5 469 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=88570 $D=1
M459 6 470 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=93200 $D=1
M460 471 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=88570 $D=1
M461 472 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=93200 $D=1
M462 469 465 471 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=88570 $D=1
M463 470 466 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=93200 $D=1
M464 471 83 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=88570 $D=1
M465 472 83 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=93200 $D=1
M466 253 84 471 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=88570 $D=1
M467 254 84 472 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=93200 $D=1
M468 473 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=88570 $D=1
M469 474 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=93200 $D=1
M470 5 85 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=88570 $D=1
M471 6 85 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=93200 $D=1
M472 477 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=88570 $D=1
M473 478 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=93200 $D=1
M474 479 85 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=88570 $D=1
M475 480 85 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=93200 $D=1
M476 5 479 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=88570 $D=1
M477 6 480 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=93200 $D=1
M478 481 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=88570 $D=1
M479 482 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=93200 $D=1
M480 479 475 481 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=88570 $D=1
M481 480 476 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=93200 $D=1
M482 481 86 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=88570 $D=1
M483 482 86 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=93200 $D=1
M484 253 87 481 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=88570 $D=1
M485 254 87 482 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=93200 $D=1
M486 483 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=88570 $D=1
M487 484 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=93200 $D=1
M488 5 88 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=88570 $D=1
M489 6 88 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=93200 $D=1
M490 487 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=88570 $D=1
M491 488 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=93200 $D=1
M492 489 88 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=88570 $D=1
M493 490 88 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=93200 $D=1
M494 5 489 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=88570 $D=1
M495 6 490 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=93200 $D=1
M496 491 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=88570 $D=1
M497 492 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=93200 $D=1
M498 489 485 491 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=88570 $D=1
M499 490 486 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=93200 $D=1
M500 491 89 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=88570 $D=1
M501 492 89 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=93200 $D=1
M502 253 90 491 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=88570 $D=1
M503 254 90 492 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=93200 $D=1
M504 493 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=88570 $D=1
M505 494 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=93200 $D=1
M506 5 91 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=88570 $D=1
M507 6 91 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=93200 $D=1
M508 497 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=88570 $D=1
M509 498 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=93200 $D=1
M510 499 91 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=88570 $D=1
M511 500 91 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=93200 $D=1
M512 5 499 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=88570 $D=1
M513 6 500 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=93200 $D=1
M514 501 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=88570 $D=1
M515 502 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=93200 $D=1
M516 499 495 501 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=88570 $D=1
M517 500 496 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=93200 $D=1
M518 501 92 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=88570 $D=1
M519 502 92 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=93200 $D=1
M520 253 93 501 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=88570 $D=1
M521 254 93 502 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=93200 $D=1
M522 503 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=88570 $D=1
M523 504 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=93200 $D=1
M524 5 94 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=88570 $D=1
M525 6 94 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=93200 $D=1
M526 507 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=88570 $D=1
M527 508 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=93200 $D=1
M528 509 94 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=88570 $D=1
M529 510 94 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=93200 $D=1
M530 5 509 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=88570 $D=1
M531 6 510 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=93200 $D=1
M532 511 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=88570 $D=1
M533 512 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=93200 $D=1
M534 509 505 511 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=88570 $D=1
M535 510 506 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=93200 $D=1
M536 511 95 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=88570 $D=1
M537 512 95 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=93200 $D=1
M538 253 96 511 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=88570 $D=1
M539 254 96 512 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=93200 $D=1
M540 513 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=88570 $D=1
M541 514 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=93200 $D=1
M542 5 97 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=88570 $D=1
M543 6 97 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=93200 $D=1
M544 517 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=88570 $D=1
M545 518 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=93200 $D=1
M546 519 97 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=88570 $D=1
M547 520 97 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=93200 $D=1
M548 5 519 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=88570 $D=1
M549 6 520 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=93200 $D=1
M550 521 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=88570 $D=1
M551 522 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=93200 $D=1
M552 519 515 521 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=88570 $D=1
M553 520 516 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=93200 $D=1
M554 521 98 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=88570 $D=1
M555 522 98 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=93200 $D=1
M556 253 99 521 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=88570 $D=1
M557 254 99 522 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=93200 $D=1
M558 523 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=88570 $D=1
M559 524 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=93200 $D=1
M560 5 100 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=88570 $D=1
M561 6 100 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=93200 $D=1
M562 527 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=88570 $D=1
M563 528 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=93200 $D=1
M564 529 100 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=88570 $D=1
M565 530 100 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=93200 $D=1
M566 5 529 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=88570 $D=1
M567 6 530 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=93200 $D=1
M568 531 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=88570 $D=1
M569 532 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=93200 $D=1
M570 529 525 531 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=88570 $D=1
M571 530 526 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=93200 $D=1
M572 531 101 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=88570 $D=1
M573 532 101 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=93200 $D=1
M574 253 102 531 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=88570 $D=1
M575 254 102 532 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=93200 $D=1
M576 533 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=88570 $D=1
M577 534 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=93200 $D=1
M578 5 103 535 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=88570 $D=1
M579 6 103 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=93200 $D=1
M580 537 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=88570 $D=1
M581 538 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=93200 $D=1
M582 539 103 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=88570 $D=1
M583 540 103 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=93200 $D=1
M584 5 539 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=88570 $D=1
M585 6 540 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=93200 $D=1
M586 541 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=88570 $D=1
M587 542 773 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=93200 $D=1
M588 539 535 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=88570 $D=1
M589 540 536 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=93200 $D=1
M590 541 104 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=88570 $D=1
M591 542 104 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=93200 $D=1
M592 253 105 541 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=88570 $D=1
M593 254 105 542 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=93200 $D=1
M594 543 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=88570 $D=1
M595 544 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=93200 $D=1
M596 5 106 545 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=88570 $D=1
M597 6 106 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=93200 $D=1
M598 547 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=88570 $D=1
M599 548 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=93200 $D=1
M600 549 106 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=88570 $D=1
M601 550 106 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=93200 $D=1
M602 5 549 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=88570 $D=1
M603 6 550 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=93200 $D=1
M604 551 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=88570 $D=1
M605 552 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=93200 $D=1
M606 549 545 551 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=88570 $D=1
M607 550 546 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=93200 $D=1
M608 551 107 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=88570 $D=1
M609 552 107 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=93200 $D=1
M610 253 108 551 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=88570 $D=1
M611 254 108 552 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=93200 $D=1
M612 553 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=88570 $D=1
M613 554 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=93200 $D=1
M614 5 109 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=88570 $D=1
M615 6 109 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=93200 $D=1
M616 557 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=88570 $D=1
M617 558 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=93200 $D=1
M618 5 110 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=88570 $D=1
M619 6 110 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=93200 $D=1
M620 253 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=88570 $D=1
M621 254 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=93200 $D=1
M622 5 561 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=88570 $D=1
M623 6 562 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=93200 $D=1
M624 561 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=88570 $D=1
M625 562 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=93200 $D=1
M626 776 249 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=88570 $D=1
M627 777 250 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=93200 $D=1
M628 563 559 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=88570 $D=1
M629 564 560 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=93200 $D=1
M630 5 563 565 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=88570 $D=1
M631 6 564 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=93200 $D=1
M632 778 565 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=88570 $D=1
M633 779 566 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=93200 $D=1
M634 563 561 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=88570 $D=1
M635 564 562 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=93200 $D=1
M636 5 569 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=88570 $D=1
M637 6 570 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=93200 $D=1
M638 569 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=88570 $D=1
M639 570 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=93200 $D=1
M640 780 253 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=88570 $D=1
M641 781 254 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=93200 $D=1
M642 571 567 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=88570 $D=1
M643 572 568 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=93200 $D=1
M644 5 571 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=88570 $D=1
M645 6 572 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=93200 $D=1
M646 782 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=88570 $D=1
M647 783 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=93200 $D=1
M648 571 569 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=88570 $D=1
M649 572 570 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=93200 $D=1
M650 573 118 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=88570 $D=1
M651 574 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=93200 $D=1
M652 575 573 565 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=88570 $D=1
M653 576 574 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=93200 $D=1
M654 119 118 575 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=88570 $D=1
M655 119 118 576 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=93200 $D=1
M656 577 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=88570 $D=1
M657 578 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=93200 $D=1
M658 579 577 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=88570 $D=1
M659 580 578 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=93200 $D=1
M660 784 120 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=88570 $D=1
M661 785 120 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=93200 $D=1
M662 5 112 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=88570 $D=1
M663 6 113 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=93200 $D=1
M664 581 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=88570 $D=1
M665 582 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=93200 $D=1
M666 583 581 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=88570 $D=1
M667 584 582 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=93200 $D=1
M668 10 122 583 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=88570 $D=1
M669 11 122 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=93200 $D=1
M670 586 585 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=88570 $D=1
M671 587 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=93200 $D=1
M672 5 590 588 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=88570 $D=1
M673 6 591 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=93200 $D=1
M674 592 575 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=88570 $D=1
M675 593 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=93200 $D=1
M676 590 592 585 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=88570 $D=1
M677 591 593 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=93200 $D=1
M678 586 575 590 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=88570 $D=1
M679 587 576 591 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=93200 $D=1
M680 594 588 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=88570 $D=1
M681 595 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=93200 $D=1
M682 596 594 583 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=88570 $D=1
M683 585 595 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=93200 $D=1
M684 575 588 596 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=88570 $D=1
M685 576 589 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=93200 $D=1
M686 597 596 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=88570 $D=1
M687 598 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=93200 $D=1
M688 599 588 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=88570 $D=1
M689 600 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=93200 $D=1
M690 601 599 597 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=88570 $D=1
M691 602 600 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=93200 $D=1
M692 583 588 601 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=88570 $D=1
M693 584 589 602 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=93200 $D=1
M694 603 575 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=88570 $D=1
M695 604 576 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=93200 $D=1
M696 5 583 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=88570 $D=1
M697 6 584 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=93200 $D=1
M698 605 601 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=88570 $D=1
M699 606 602 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=93200 $D=1
M700 804 575 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=88570 $D=1
M701 805 576 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=93200 $D=1
M702 607 583 804 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=88570 $D=1
M703 608 584 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=93200 $D=1
M704 806 575 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=88570 $D=1
M705 807 576 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=93200 $D=1
M706 609 583 806 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=88570 $D=1
M707 610 584 807 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=93200 $D=1
M708 613 575 611 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=88570 $D=1
M709 614 576 612 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=93200 $D=1
M710 611 583 613 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=88570 $D=1
M711 612 584 614 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=93200 $D=1
M712 5 609 611 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=88570 $D=1
M713 6 610 612 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=93200 $D=1
M714 615 126 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=88570 $D=1
M715 616 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=93200 $D=1
M716 617 615 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=88570 $D=1
M717 618 616 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=93200 $D=1
M718 607 126 617 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=88570 $D=1
M719 608 126 618 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=93200 $D=1
M720 619 615 605 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=88570 $D=1
M721 620 616 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=93200 $D=1
M722 613 126 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=88570 $D=1
M723 614 126 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=93200 $D=1
M724 621 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=88570 $D=1
M725 622 127 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=93200 $D=1
M726 623 621 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=88570 $D=1
M727 624 622 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=93200 $D=1
M728 617 127 623 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=88570 $D=1
M729 618 127 624 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=93200 $D=1
M730 12 623 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=88570 $D=1
M731 13 624 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=93200 $D=1
M732 625 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=88570 $D=1
M733 626 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=93200 $D=1
M734 627 625 129 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=88570 $D=1
M735 628 626 130 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=93200 $D=1
M736 131 128 627 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=88570 $D=1
M737 132 128 628 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=93200 $D=1
M738 629 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=88570 $D=1
M739 630 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=93200 $D=1
M740 631 629 133 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=88570 $D=1
M741 632 630 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=93200 $D=1
M742 135 128 631 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=88570 $D=1
M743 136 128 632 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=93200 $D=1
M744 633 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=88570 $D=1
M745 634 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=93200 $D=1
M746 635 633 136 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=88570 $D=1
M747 636 634 137 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=93200 $D=1
M748 114 128 635 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=88570 $D=1
M749 116 128 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=93200 $D=1
M750 637 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=88570 $D=1
M751 638 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=93200 $D=1
M752 639 637 138 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=88570 $D=1
M753 640 638 139 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=93200 $D=1
M754 115 128 639 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=88570 $D=1
M755 117 128 640 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=93200 $D=1
M756 641 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=88570 $D=1
M757 642 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=93200 $D=1
M758 643 641 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=88570 $D=1
M759 644 642 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=93200 $D=1
M760 140 128 643 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=88570 $D=1
M761 141 128 644 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=93200 $D=1
M762 5 575 786 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=88570 $D=1
M763 6 576 787 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=93200 $D=1
M764 132 786 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=88570 $D=1
M765 129 787 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=93200 $D=1
M766 645 142 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=88570 $D=1
M767 646 142 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=93200 $D=1
M768 143 645 132 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=88570 $D=1
M769 144 646 129 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=93200 $D=1
M770 627 142 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=88570 $D=1
M771 628 142 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=93200 $D=1
M772 647 145 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=88570 $D=1
M773 648 145 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=93200 $D=1
M774 121 647 143 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=88570 $D=1
M775 146 648 144 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=93200 $D=1
M776 631 145 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=88570 $D=1
M777 632 145 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=93200 $D=1
M778 649 147 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=88570 $D=1
M779 650 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=93200 $D=1
M780 124 649 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=88570 $D=1
M781 125 650 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=93200 $D=1
M782 635 147 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=88570 $D=1
M783 636 147 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=93200 $D=1
M784 651 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=88570 $D=1
M785 652 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=93200 $D=1
M786 149 651 124 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=88570 $D=1
M787 150 652 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=93200 $D=1
M788 639 148 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=88570 $D=1
M789 640 148 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=93200 $D=1
M790 653 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=88570 $D=1
M791 654 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=93200 $D=1
M792 225 653 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=88570 $D=1
M793 226 654 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=93200 $D=1
M794 643 151 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=88570 $D=1
M795 644 151 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=93200 $D=1
M796 655 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=88570 $D=1
M797 656 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=93200 $D=1
M798 657 655 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=88570 $D=1
M799 658 656 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=93200 $D=1
M800 10 152 657 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=88570 $D=1
M801 11 152 658 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=93200 $D=1
M802 808 565 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=88570 $D=1
M803 809 566 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=93200 $D=1
M804 659 657 808 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=88570 $D=1
M805 660 658 809 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=93200 $D=1
M806 663 565 661 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=88570 $D=1
M807 664 566 662 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=93200 $D=1
M808 661 657 663 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=88570 $D=1
M809 662 658 664 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=93200 $D=1
M810 5 659 661 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=88570 $D=1
M811 6 660 662 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=93200 $D=1
M812 810 153 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=88570 $D=1
M813 811 665 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=93200 $D=1
M814 788 663 810 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=88570 $D=1
M815 789 664 811 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=93200 $D=1
M816 665 788 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=88570 $D=1
M817 154 789 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=93200 $D=1
M818 666 565 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=88570 $D=1
M819 667 566 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=93200 $D=1
M820 5 668 666 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=88570 $D=1
M821 6 669 667 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=93200 $D=1
M822 668 657 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=88570 $D=1
M823 669 658 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=93200 $D=1
M824 812 666 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=88570 $D=1
M825 813 667 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=93200 $D=1
M826 670 153 812 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=88570 $D=1
M827 671 665 813 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=93200 $D=1
M828 673 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=88570 $D=1
M829 674 672 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=93200 $D=1
M830 814 670 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=88570 $D=1
M831 815 671 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=93200 $D=1
M832 672 673 814 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=88570 $D=1
M833 156 674 815 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=93200 $D=1
M834 676 675 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=88570 $D=1
M835 677 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=93200 $D=1
M836 5 680 678 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=88570 $D=1
M837 6 681 679 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=93200 $D=1
M838 682 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=88570 $D=1
M839 683 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=93200 $D=1
M840 680 682 675 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=88570 $D=1
M841 681 683 157 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=93200 $D=1
M842 676 119 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=88570 $D=1
M843 677 119 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=93200 $D=1
M844 684 678 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=88570 $D=1
M845 685 679 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=93200 $D=1
M846 158 684 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=88570 $D=1
M847 675 685 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=93200 $D=1
M848 119 678 158 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=88570 $D=1
M849 119 679 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=93200 $D=1
M850 686 158 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=88570 $D=1
M851 687 675 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=93200 $D=1
M852 688 678 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=88570 $D=1
M853 689 679 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=93200 $D=1
M854 227 688 686 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=88570 $D=1
M855 228 689 687 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=93200 $D=1
M856 5 678 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=88570 $D=1
M857 6 679 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=93200 $D=1
M858 690 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=88570 $D=1
M859 691 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=93200 $D=1
M860 692 690 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=88570 $D=1
M861 693 691 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=93200 $D=1
M862 12 159 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=88570 $D=1
M863 13 159 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=93200 $D=1
M864 694 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=88570 $D=1
M865 695 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=93200 $D=1
M866 160 694 692 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=88570 $D=1
M867 160 695 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=93200 $D=1
M868 5 160 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=88570 $D=1
M869 6 160 160 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=93200 $D=1
M870 696 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=88570 $D=1
M871 697 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=93200 $D=1
M872 5 696 698 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=88570 $D=1
M873 6 697 699 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=93200 $D=1
M874 700 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=88570 $D=1
M875 701 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=93200 $D=1
M876 702 696 160 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=88570 $D=1
M877 703 697 160 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=93200 $D=1
M878 5 702 790 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=88570 $D=1
M879 6 703 791 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=93200 $D=1
M880 704 790 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=88570 $D=1
M881 705 791 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=93200 $D=1
M882 702 698 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=88570 $D=1
M883 703 699 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=93200 $D=1
M884 706 111 704 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=88570 $D=1
M885 707 111 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=93200 $D=1
M886 5 710 708 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=88570 $D=1
M887 6 711 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=93200 $D=1
M888 710 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=88570 $D=1
M889 711 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=93200 $D=1
M890 792 706 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=88570 $D=1
M891 793 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=93200 $D=1
M892 712 708 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=88570 $D=1
M893 713 709 793 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=93200 $D=1
M894 5 712 119 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=88570 $D=1
M895 6 713 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=93200 $D=1
M896 794 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=88570 $D=1
M897 795 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=93200 $D=1
M898 712 710 794 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=88570 $D=1
M899 713 711 795 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=93200 $D=1
M900 201 1 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=89820 $D=0
M901 202 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=94450 $D=0
M902 203 1 2 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=89820 $D=0
M903 204 1 3 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=94450 $D=0
M904 5 201 203 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=89820 $D=0
M905 6 202 204 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=94450 $D=0
M906 205 1 4 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=89820 $D=0
M907 206 1 4 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=94450 $D=0
M908 2 201 205 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=89820 $D=0
M909 3 202 206 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=94450 $D=0
M910 207 1 5 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=89820 $D=0
M911 208 1 6 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=94450 $D=0
M912 2 201 207 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=89820 $D=0
M913 3 202 208 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=94450 $D=0
M914 211 7 207 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=89820 $D=0
M915 212 7 208 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=94450 $D=0
M916 209 7 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=89820 $D=0
M917 210 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=94450 $D=0
M918 213 7 205 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=89820 $D=0
M919 214 7 206 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=94450 $D=0
M920 203 209 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=89820 $D=0
M921 204 210 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=94450 $D=0
M922 215 8 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=89820 $D=0
M923 216 8 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=94450 $D=0
M924 217 8 213 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=89820 $D=0
M925 218 8 214 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=94450 $D=0
M926 211 215 217 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=89820 $D=0
M927 212 216 218 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=94450 $D=0
M928 219 9 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=89820 $D=0
M929 220 9 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=94450 $D=0
M930 221 9 5 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=89820 $D=0
M931 222 9 6 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=94450 $D=0
M932 10 219 221 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=89820 $D=0
M933 11 220 222 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=94450 $D=0
M934 223 9 12 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=89820 $D=0
M935 224 9 13 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=94450 $D=0
M936 225 219 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=89820 $D=0
M937 226 220 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=94450 $D=0
M938 229 9 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=89820 $D=0
M939 230 9 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=94450 $D=0
M940 217 219 229 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=89820 $D=0
M941 218 220 230 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=94450 $D=0
M942 233 14 229 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=89820 $D=0
M943 234 14 230 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=94450 $D=0
M944 231 14 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=89820 $D=0
M945 232 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=94450 $D=0
M946 235 14 223 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=89820 $D=0
M947 236 14 224 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=94450 $D=0
M948 221 231 235 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=89820 $D=0
M949 222 232 236 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=94450 $D=0
M950 237 15 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=89820 $D=0
M951 238 15 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=94450 $D=0
M952 239 15 235 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=89820 $D=0
M953 240 15 236 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=94450 $D=0
M954 233 237 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=89820 $D=0
M955 234 238 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=94450 $D=0
M956 161 16 241 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=89820 $D=0
M957 162 16 242 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=94450 $D=0
M958 243 17 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=89820 $D=0
M959 244 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=94450 $D=0
M960 245 241 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=89820 $D=0
M961 246 242 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=94450 $D=0
M962 161 245 714 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=89820 $D=0
M963 162 246 715 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=94450 $D=0
M964 247 714 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=89820 $D=0
M965 248 715 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=94450 $D=0
M966 245 16 247 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=89820 $D=0
M967 246 16 248 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=94450 $D=0
M968 247 243 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=89820 $D=0
M969 248 244 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=94450 $D=0
M970 253 251 247 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=89820 $D=0
M971 254 252 248 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=94450 $D=0
M972 251 18 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=89820 $D=0
M973 252 18 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=94450 $D=0
M974 161 19 255 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=89820 $D=0
M975 162 19 256 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=94450 $D=0
M976 257 20 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=89820 $D=0
M977 258 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=94450 $D=0
M978 259 255 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=89820 $D=0
M979 260 256 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=94450 $D=0
M980 161 259 716 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=89820 $D=0
M981 162 260 717 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=94450 $D=0
M982 261 716 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=89820 $D=0
M983 262 717 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=94450 $D=0
M984 259 19 261 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=89820 $D=0
M985 260 19 262 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=94450 $D=0
M986 261 257 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=89820 $D=0
M987 262 258 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=94450 $D=0
M988 253 263 261 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=89820 $D=0
M989 254 264 262 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=94450 $D=0
M990 263 21 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=89820 $D=0
M991 264 21 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=94450 $D=0
M992 161 22 265 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=89820 $D=0
M993 162 22 266 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=94450 $D=0
M994 267 23 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=89820 $D=0
M995 268 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=94450 $D=0
M996 269 265 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=89820 $D=0
M997 270 266 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=94450 $D=0
M998 161 269 718 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=89820 $D=0
M999 162 270 719 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=94450 $D=0
M1000 271 718 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=89820 $D=0
M1001 272 719 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=94450 $D=0
M1002 269 22 271 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=89820 $D=0
M1003 270 22 272 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=94450 $D=0
M1004 271 267 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=89820 $D=0
M1005 272 268 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=94450 $D=0
M1006 253 273 271 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=89820 $D=0
M1007 254 274 272 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=94450 $D=0
M1008 273 24 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=89820 $D=0
M1009 274 24 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=94450 $D=0
M1010 161 25 275 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=89820 $D=0
M1011 162 25 276 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=94450 $D=0
M1012 277 26 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=89820 $D=0
M1013 278 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=94450 $D=0
M1014 279 275 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=89820 $D=0
M1015 280 276 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=94450 $D=0
M1016 161 279 720 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=89820 $D=0
M1017 162 280 721 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=94450 $D=0
M1018 281 720 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=89820 $D=0
M1019 282 721 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=94450 $D=0
M1020 279 25 281 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=89820 $D=0
M1021 280 25 282 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=94450 $D=0
M1022 281 277 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=89820 $D=0
M1023 282 278 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=94450 $D=0
M1024 253 283 281 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=89820 $D=0
M1025 254 284 282 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=94450 $D=0
M1026 283 27 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=89820 $D=0
M1027 284 27 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=94450 $D=0
M1028 161 28 285 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=89820 $D=0
M1029 162 28 286 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=94450 $D=0
M1030 287 29 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=89820 $D=0
M1031 288 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=94450 $D=0
M1032 289 285 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=89820 $D=0
M1033 290 286 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=94450 $D=0
M1034 161 289 722 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=89820 $D=0
M1035 162 290 723 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=94450 $D=0
M1036 291 722 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=89820 $D=0
M1037 292 723 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=94450 $D=0
M1038 289 28 291 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=89820 $D=0
M1039 290 28 292 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=94450 $D=0
M1040 291 287 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=89820 $D=0
M1041 292 288 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=94450 $D=0
M1042 253 293 291 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=89820 $D=0
M1043 254 294 292 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=94450 $D=0
M1044 293 30 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=89820 $D=0
M1045 294 30 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=94450 $D=0
M1046 161 31 295 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=89820 $D=0
M1047 162 31 296 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=94450 $D=0
M1048 297 32 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=89820 $D=0
M1049 298 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=94450 $D=0
M1050 299 295 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=89820 $D=0
M1051 300 296 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=94450 $D=0
M1052 161 299 724 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=89820 $D=0
M1053 162 300 725 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=94450 $D=0
M1054 301 724 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=89820 $D=0
M1055 302 725 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=94450 $D=0
M1056 299 31 301 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=89820 $D=0
M1057 300 31 302 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=94450 $D=0
M1058 301 297 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=89820 $D=0
M1059 302 298 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=94450 $D=0
M1060 253 303 301 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=89820 $D=0
M1061 254 304 302 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=94450 $D=0
M1062 303 33 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=89820 $D=0
M1063 304 33 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=94450 $D=0
M1064 161 34 305 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=89820 $D=0
M1065 162 34 306 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=94450 $D=0
M1066 307 35 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=89820 $D=0
M1067 308 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=94450 $D=0
M1068 309 305 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=89820 $D=0
M1069 310 306 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=94450 $D=0
M1070 161 309 726 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=89820 $D=0
M1071 162 310 727 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=94450 $D=0
M1072 311 726 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=89820 $D=0
M1073 312 727 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=94450 $D=0
M1074 309 34 311 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=89820 $D=0
M1075 310 34 312 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=94450 $D=0
M1076 311 307 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=89820 $D=0
M1077 312 308 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=94450 $D=0
M1078 253 313 311 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=89820 $D=0
M1079 254 314 312 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=94450 $D=0
M1080 313 36 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=89820 $D=0
M1081 314 36 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=94450 $D=0
M1082 161 37 315 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=89820 $D=0
M1083 162 37 316 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=94450 $D=0
M1084 317 38 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=89820 $D=0
M1085 318 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=94450 $D=0
M1086 319 315 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=89820 $D=0
M1087 320 316 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=94450 $D=0
M1088 161 319 728 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=89820 $D=0
M1089 162 320 729 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=94450 $D=0
M1090 321 728 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=89820 $D=0
M1091 322 729 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=94450 $D=0
M1092 319 37 321 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=89820 $D=0
M1093 320 37 322 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=94450 $D=0
M1094 321 317 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=89820 $D=0
M1095 322 318 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=94450 $D=0
M1096 253 323 321 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=89820 $D=0
M1097 254 324 322 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=94450 $D=0
M1098 323 39 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=89820 $D=0
M1099 324 39 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=94450 $D=0
M1100 161 40 325 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=89820 $D=0
M1101 162 40 326 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=94450 $D=0
M1102 327 41 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=89820 $D=0
M1103 328 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=94450 $D=0
M1104 329 325 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=89820 $D=0
M1105 330 326 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=94450 $D=0
M1106 161 329 730 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=89820 $D=0
M1107 162 330 731 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=94450 $D=0
M1108 331 730 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=89820 $D=0
M1109 332 731 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=94450 $D=0
M1110 329 40 331 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=89820 $D=0
M1111 330 40 332 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=94450 $D=0
M1112 331 327 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=89820 $D=0
M1113 332 328 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=94450 $D=0
M1114 253 333 331 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=89820 $D=0
M1115 254 334 332 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=94450 $D=0
M1116 333 42 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=89820 $D=0
M1117 334 42 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=94450 $D=0
M1118 161 43 335 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=89820 $D=0
M1119 162 43 336 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=94450 $D=0
M1120 337 44 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=89820 $D=0
M1121 338 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=94450 $D=0
M1122 339 335 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=89820 $D=0
M1123 340 336 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=94450 $D=0
M1124 161 339 732 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=89820 $D=0
M1125 162 340 733 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=94450 $D=0
M1126 341 732 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=89820 $D=0
M1127 342 733 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=94450 $D=0
M1128 339 43 341 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=89820 $D=0
M1129 340 43 342 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=94450 $D=0
M1130 341 337 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=89820 $D=0
M1131 342 338 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=94450 $D=0
M1132 253 343 341 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=89820 $D=0
M1133 254 344 342 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=94450 $D=0
M1134 343 45 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=89820 $D=0
M1135 344 45 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=94450 $D=0
M1136 161 46 345 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=89820 $D=0
M1137 162 46 346 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=94450 $D=0
M1138 347 47 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=89820 $D=0
M1139 348 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=94450 $D=0
M1140 349 345 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=89820 $D=0
M1141 350 346 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=94450 $D=0
M1142 161 349 734 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=89820 $D=0
M1143 162 350 735 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=94450 $D=0
M1144 351 734 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=89820 $D=0
M1145 352 735 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=94450 $D=0
M1146 349 46 351 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=89820 $D=0
M1147 350 46 352 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=94450 $D=0
M1148 351 347 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=89820 $D=0
M1149 352 348 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=94450 $D=0
M1150 253 353 351 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=89820 $D=0
M1151 254 354 352 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=94450 $D=0
M1152 353 48 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=89820 $D=0
M1153 354 48 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=94450 $D=0
M1154 161 49 355 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=89820 $D=0
M1155 162 49 356 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=94450 $D=0
M1156 357 50 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=89820 $D=0
M1157 358 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=94450 $D=0
M1158 359 355 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=89820 $D=0
M1159 360 356 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=94450 $D=0
M1160 161 359 736 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=89820 $D=0
M1161 162 360 737 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=94450 $D=0
M1162 361 736 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=89820 $D=0
M1163 362 737 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=94450 $D=0
M1164 359 49 361 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=89820 $D=0
M1165 360 49 362 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=94450 $D=0
M1166 361 357 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=89820 $D=0
M1167 362 358 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=94450 $D=0
M1168 253 363 361 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=89820 $D=0
M1169 254 364 362 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=94450 $D=0
M1170 363 51 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=89820 $D=0
M1171 364 51 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=94450 $D=0
M1172 161 52 365 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=89820 $D=0
M1173 162 52 366 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=94450 $D=0
M1174 367 53 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=89820 $D=0
M1175 368 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=94450 $D=0
M1176 369 365 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=89820 $D=0
M1177 370 366 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=94450 $D=0
M1178 161 369 738 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=89820 $D=0
M1179 162 370 739 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=94450 $D=0
M1180 371 738 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=89820 $D=0
M1181 372 739 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=94450 $D=0
M1182 369 52 371 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=89820 $D=0
M1183 370 52 372 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=94450 $D=0
M1184 371 367 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=89820 $D=0
M1185 372 368 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=94450 $D=0
M1186 253 373 371 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=89820 $D=0
M1187 254 374 372 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=94450 $D=0
M1188 373 54 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=89820 $D=0
M1189 374 54 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=94450 $D=0
M1190 161 55 375 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=89820 $D=0
M1191 162 55 376 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=94450 $D=0
M1192 377 56 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=89820 $D=0
M1193 378 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=94450 $D=0
M1194 379 375 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=89820 $D=0
M1195 380 376 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=94450 $D=0
M1196 161 379 740 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=89820 $D=0
M1197 162 380 741 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=94450 $D=0
M1198 381 740 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=89820 $D=0
M1199 382 741 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=94450 $D=0
M1200 379 55 381 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=89820 $D=0
M1201 380 55 382 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=94450 $D=0
M1202 381 377 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=89820 $D=0
M1203 382 378 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=94450 $D=0
M1204 253 383 381 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=89820 $D=0
M1205 254 384 382 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=94450 $D=0
M1206 383 57 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=89820 $D=0
M1207 384 57 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=94450 $D=0
M1208 161 58 385 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=89820 $D=0
M1209 162 58 386 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=94450 $D=0
M1210 387 59 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=89820 $D=0
M1211 388 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=94450 $D=0
M1212 389 385 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=89820 $D=0
M1213 390 386 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=94450 $D=0
M1214 161 389 742 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=89820 $D=0
M1215 162 390 743 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=94450 $D=0
M1216 391 742 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=89820 $D=0
M1217 392 743 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=94450 $D=0
M1218 389 58 391 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=89820 $D=0
M1219 390 58 392 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=94450 $D=0
M1220 391 387 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=89820 $D=0
M1221 392 388 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=94450 $D=0
M1222 253 393 391 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=89820 $D=0
M1223 254 394 392 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=94450 $D=0
M1224 393 60 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=89820 $D=0
M1225 394 60 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=94450 $D=0
M1226 161 61 395 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=89820 $D=0
M1227 162 61 396 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=94450 $D=0
M1228 397 62 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=89820 $D=0
M1229 398 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=94450 $D=0
M1230 399 395 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=89820 $D=0
M1231 400 396 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=94450 $D=0
M1232 161 399 744 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=89820 $D=0
M1233 162 400 745 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=94450 $D=0
M1234 401 744 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=89820 $D=0
M1235 402 745 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=94450 $D=0
M1236 399 61 401 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=89820 $D=0
M1237 400 61 402 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=94450 $D=0
M1238 401 397 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=89820 $D=0
M1239 402 398 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=94450 $D=0
M1240 253 403 401 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=89820 $D=0
M1241 254 404 402 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=94450 $D=0
M1242 403 63 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=89820 $D=0
M1243 404 63 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=94450 $D=0
M1244 161 64 405 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=89820 $D=0
M1245 162 64 406 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=94450 $D=0
M1246 407 65 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=89820 $D=0
M1247 408 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=94450 $D=0
M1248 409 405 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=89820 $D=0
M1249 410 406 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=94450 $D=0
M1250 161 409 746 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=89820 $D=0
M1251 162 410 747 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=94450 $D=0
M1252 411 746 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=89820 $D=0
M1253 412 747 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=94450 $D=0
M1254 409 64 411 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=89820 $D=0
M1255 410 64 412 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=94450 $D=0
M1256 411 407 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=89820 $D=0
M1257 412 408 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=94450 $D=0
M1258 253 413 411 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=89820 $D=0
M1259 254 414 412 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=94450 $D=0
M1260 413 66 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=89820 $D=0
M1261 414 66 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=94450 $D=0
M1262 161 67 415 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=89820 $D=0
M1263 162 67 416 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=94450 $D=0
M1264 417 68 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=89820 $D=0
M1265 418 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=94450 $D=0
M1266 419 415 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=89820 $D=0
M1267 420 416 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=94450 $D=0
M1268 161 419 748 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=89820 $D=0
M1269 162 420 749 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=94450 $D=0
M1270 421 748 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=89820 $D=0
M1271 422 749 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=94450 $D=0
M1272 419 67 421 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=89820 $D=0
M1273 420 67 422 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=94450 $D=0
M1274 421 417 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=89820 $D=0
M1275 422 418 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=94450 $D=0
M1276 253 423 421 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=89820 $D=0
M1277 254 424 422 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=94450 $D=0
M1278 423 69 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=89820 $D=0
M1279 424 69 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=94450 $D=0
M1280 161 70 425 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=89820 $D=0
M1281 162 70 426 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=94450 $D=0
M1282 427 71 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=89820 $D=0
M1283 428 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=94450 $D=0
M1284 429 425 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=89820 $D=0
M1285 430 426 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=94450 $D=0
M1286 161 429 750 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=89820 $D=0
M1287 162 430 751 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=94450 $D=0
M1288 431 750 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=89820 $D=0
M1289 432 751 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=94450 $D=0
M1290 429 70 431 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=89820 $D=0
M1291 430 70 432 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=94450 $D=0
M1292 431 427 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=89820 $D=0
M1293 432 428 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=94450 $D=0
M1294 253 433 431 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=89820 $D=0
M1295 254 434 432 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=94450 $D=0
M1296 433 72 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=89820 $D=0
M1297 434 72 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=94450 $D=0
M1298 161 73 435 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=89820 $D=0
M1299 162 73 436 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=94450 $D=0
M1300 437 74 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=89820 $D=0
M1301 438 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=94450 $D=0
M1302 439 435 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=89820 $D=0
M1303 440 436 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=94450 $D=0
M1304 161 439 752 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=89820 $D=0
M1305 162 440 753 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=94450 $D=0
M1306 441 752 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=89820 $D=0
M1307 442 753 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=94450 $D=0
M1308 439 73 441 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=89820 $D=0
M1309 440 73 442 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=94450 $D=0
M1310 441 437 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=89820 $D=0
M1311 442 438 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=94450 $D=0
M1312 253 443 441 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=89820 $D=0
M1313 254 444 442 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=94450 $D=0
M1314 443 75 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=89820 $D=0
M1315 444 75 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=94450 $D=0
M1316 161 76 445 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=89820 $D=0
M1317 162 76 446 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=94450 $D=0
M1318 447 77 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=89820 $D=0
M1319 448 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=94450 $D=0
M1320 449 445 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=89820 $D=0
M1321 450 446 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=94450 $D=0
M1322 161 449 754 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=89820 $D=0
M1323 162 450 755 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=94450 $D=0
M1324 451 754 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=89820 $D=0
M1325 452 755 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=94450 $D=0
M1326 449 76 451 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=89820 $D=0
M1327 450 76 452 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=94450 $D=0
M1328 451 447 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=89820 $D=0
M1329 452 448 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=94450 $D=0
M1330 253 453 451 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=89820 $D=0
M1331 254 454 452 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=94450 $D=0
M1332 453 78 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=89820 $D=0
M1333 454 78 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=94450 $D=0
M1334 161 79 455 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=89820 $D=0
M1335 162 79 456 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=94450 $D=0
M1336 457 80 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=89820 $D=0
M1337 458 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=94450 $D=0
M1338 459 455 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=89820 $D=0
M1339 460 456 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=94450 $D=0
M1340 161 459 756 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=89820 $D=0
M1341 162 460 757 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=94450 $D=0
M1342 461 756 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=89820 $D=0
M1343 462 757 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=94450 $D=0
M1344 459 79 461 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=89820 $D=0
M1345 460 79 462 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=94450 $D=0
M1346 461 457 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=89820 $D=0
M1347 462 458 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=94450 $D=0
M1348 253 463 461 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=89820 $D=0
M1349 254 464 462 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=94450 $D=0
M1350 463 81 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=89820 $D=0
M1351 464 81 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=94450 $D=0
M1352 161 82 465 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=89820 $D=0
M1353 162 82 466 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=94450 $D=0
M1354 467 83 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=89820 $D=0
M1355 468 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=94450 $D=0
M1356 469 465 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=89820 $D=0
M1357 470 466 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=94450 $D=0
M1358 161 469 758 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=89820 $D=0
M1359 162 470 759 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=94450 $D=0
M1360 471 758 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=89820 $D=0
M1361 472 759 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=94450 $D=0
M1362 469 82 471 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=89820 $D=0
M1363 470 82 472 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=94450 $D=0
M1364 471 467 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=89820 $D=0
M1365 472 468 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=94450 $D=0
M1366 253 473 471 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=89820 $D=0
M1367 254 474 472 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=94450 $D=0
M1368 473 84 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=89820 $D=0
M1369 474 84 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=94450 $D=0
M1370 161 85 475 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=89820 $D=0
M1371 162 85 476 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=94450 $D=0
M1372 477 86 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=89820 $D=0
M1373 478 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=94450 $D=0
M1374 479 475 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=89820 $D=0
M1375 480 476 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=94450 $D=0
M1376 161 479 760 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=89820 $D=0
M1377 162 480 761 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=94450 $D=0
M1378 481 760 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=89820 $D=0
M1379 482 761 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=94450 $D=0
M1380 479 85 481 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=89820 $D=0
M1381 480 85 482 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=94450 $D=0
M1382 481 477 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=89820 $D=0
M1383 482 478 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=94450 $D=0
M1384 253 483 481 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=89820 $D=0
M1385 254 484 482 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=94450 $D=0
M1386 483 87 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=89820 $D=0
M1387 484 87 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=94450 $D=0
M1388 161 88 485 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=89820 $D=0
M1389 162 88 486 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=94450 $D=0
M1390 487 89 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=89820 $D=0
M1391 488 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=94450 $D=0
M1392 489 485 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=89820 $D=0
M1393 490 486 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=94450 $D=0
M1394 161 489 762 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=89820 $D=0
M1395 162 490 763 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=94450 $D=0
M1396 491 762 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=89820 $D=0
M1397 492 763 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=94450 $D=0
M1398 489 88 491 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=89820 $D=0
M1399 490 88 492 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=94450 $D=0
M1400 491 487 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=89820 $D=0
M1401 492 488 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=94450 $D=0
M1402 253 493 491 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=89820 $D=0
M1403 254 494 492 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=94450 $D=0
M1404 493 90 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=89820 $D=0
M1405 494 90 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=94450 $D=0
M1406 161 91 495 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=89820 $D=0
M1407 162 91 496 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=94450 $D=0
M1408 497 92 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=89820 $D=0
M1409 498 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=94450 $D=0
M1410 499 495 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=89820 $D=0
M1411 500 496 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=94450 $D=0
M1412 161 499 764 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=89820 $D=0
M1413 162 500 765 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=94450 $D=0
M1414 501 764 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=89820 $D=0
M1415 502 765 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=94450 $D=0
M1416 499 91 501 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=89820 $D=0
M1417 500 91 502 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=94450 $D=0
M1418 501 497 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=89820 $D=0
M1419 502 498 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=94450 $D=0
M1420 253 503 501 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=89820 $D=0
M1421 254 504 502 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=94450 $D=0
M1422 503 93 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=89820 $D=0
M1423 504 93 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=94450 $D=0
M1424 161 94 505 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=89820 $D=0
M1425 162 94 506 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=94450 $D=0
M1426 507 95 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=89820 $D=0
M1427 508 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=94450 $D=0
M1428 509 505 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=89820 $D=0
M1429 510 506 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=94450 $D=0
M1430 161 509 766 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=89820 $D=0
M1431 162 510 767 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=94450 $D=0
M1432 511 766 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=89820 $D=0
M1433 512 767 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=94450 $D=0
M1434 509 94 511 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=89820 $D=0
M1435 510 94 512 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=94450 $D=0
M1436 511 507 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=89820 $D=0
M1437 512 508 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=94450 $D=0
M1438 253 513 511 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=89820 $D=0
M1439 254 514 512 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=94450 $D=0
M1440 513 96 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=89820 $D=0
M1441 514 96 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=94450 $D=0
M1442 161 97 515 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=89820 $D=0
M1443 162 97 516 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=94450 $D=0
M1444 517 98 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=89820 $D=0
M1445 518 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=94450 $D=0
M1446 519 515 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=89820 $D=0
M1447 520 516 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=94450 $D=0
M1448 161 519 768 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=89820 $D=0
M1449 162 520 769 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=94450 $D=0
M1450 521 768 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=89820 $D=0
M1451 522 769 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=94450 $D=0
M1452 519 97 521 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=89820 $D=0
M1453 520 97 522 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=94450 $D=0
M1454 521 517 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=89820 $D=0
M1455 522 518 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=94450 $D=0
M1456 253 523 521 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=89820 $D=0
M1457 254 524 522 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=94450 $D=0
M1458 523 99 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=89820 $D=0
M1459 524 99 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=94450 $D=0
M1460 161 100 525 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=89820 $D=0
M1461 162 100 526 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=94450 $D=0
M1462 527 101 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=89820 $D=0
M1463 528 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=94450 $D=0
M1464 529 525 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=89820 $D=0
M1465 530 526 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=94450 $D=0
M1466 161 529 770 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=89820 $D=0
M1467 162 530 771 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=94450 $D=0
M1468 531 770 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=89820 $D=0
M1469 532 771 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=94450 $D=0
M1470 529 100 531 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=89820 $D=0
M1471 530 100 532 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=94450 $D=0
M1472 531 527 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=89820 $D=0
M1473 532 528 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=94450 $D=0
M1474 253 533 531 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=89820 $D=0
M1475 254 534 532 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=94450 $D=0
M1476 533 102 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=89820 $D=0
M1477 534 102 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=94450 $D=0
M1478 161 103 535 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=89820 $D=0
M1479 162 103 536 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=94450 $D=0
M1480 537 104 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=89820 $D=0
M1481 538 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=94450 $D=0
M1482 539 535 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=89820 $D=0
M1483 540 536 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=94450 $D=0
M1484 161 539 772 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=89820 $D=0
M1485 162 540 773 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=94450 $D=0
M1486 541 772 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=89820 $D=0
M1487 542 773 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=94450 $D=0
M1488 539 103 541 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=89820 $D=0
M1489 540 103 542 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=94450 $D=0
M1490 541 537 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=89820 $D=0
M1491 542 538 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=94450 $D=0
M1492 253 543 541 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=89820 $D=0
M1493 254 544 542 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=94450 $D=0
M1494 543 105 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=89820 $D=0
M1495 544 105 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=94450 $D=0
M1496 161 106 545 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=89820 $D=0
M1497 162 106 546 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=94450 $D=0
M1498 547 107 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=89820 $D=0
M1499 548 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=94450 $D=0
M1500 549 545 239 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=89820 $D=0
M1501 550 546 240 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=94450 $D=0
M1502 161 549 774 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=89820 $D=0
M1503 162 550 775 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=94450 $D=0
M1504 551 774 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=89820 $D=0
M1505 552 775 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=94450 $D=0
M1506 549 106 551 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=89820 $D=0
M1507 550 106 552 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=94450 $D=0
M1508 551 547 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=89820 $D=0
M1509 552 548 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=94450 $D=0
M1510 253 553 551 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=89820 $D=0
M1511 254 554 552 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=94450 $D=0
M1512 553 108 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=89820 $D=0
M1513 554 108 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=94450 $D=0
M1514 161 109 555 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=89820 $D=0
M1515 162 109 556 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=94450 $D=0
M1516 557 110 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=89820 $D=0
M1517 558 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=94450 $D=0
M1518 5 557 249 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=89820 $D=0
M1519 6 558 250 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=94450 $D=0
M1520 253 555 5 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=89820 $D=0
M1521 254 556 6 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=94450 $D=0
M1522 161 561 559 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=89820 $D=0
M1523 162 562 560 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=94450 $D=0
M1524 561 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=89820 $D=0
M1525 562 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=94450 $D=0
M1526 776 249 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=89820 $D=0
M1527 777 250 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=94450 $D=0
M1528 563 561 776 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=89820 $D=0
M1529 564 562 777 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=94450 $D=0
M1530 161 563 565 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=89820 $D=0
M1531 162 564 566 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=94450 $D=0
M1532 778 565 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=89820 $D=0
M1533 779 566 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=94450 $D=0
M1534 563 559 778 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=89820 $D=0
M1535 564 560 779 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=94450 $D=0
M1536 161 569 567 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=89820 $D=0
M1537 162 570 568 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=94450 $D=0
M1538 569 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=89820 $D=0
M1539 570 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=94450 $D=0
M1540 780 253 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=89820 $D=0
M1541 781 254 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=94450 $D=0
M1542 571 569 780 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=89820 $D=0
M1543 572 570 781 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=94450 $D=0
M1544 161 571 112 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=89820 $D=0
M1545 162 572 113 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=94450 $D=0
M1546 782 112 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=89820 $D=0
M1547 783 113 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=94450 $D=0
M1548 571 567 782 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=89820 $D=0
M1549 572 568 783 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=94450 $D=0
M1550 573 118 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=89820 $D=0
M1551 574 118 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=94450 $D=0
M1552 575 118 565 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=89820 $D=0
M1553 576 118 566 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=94450 $D=0
M1554 119 573 575 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=89820 $D=0
M1555 119 574 576 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=94450 $D=0
M1556 577 120 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=89820 $D=0
M1557 578 120 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=94450 $D=0
M1558 579 120 112 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=89820 $D=0
M1559 580 120 113 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=94450 $D=0
M1560 784 577 579 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=89820 $D=0
M1561 785 578 580 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=94450 $D=0
M1562 161 112 784 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=89820 $D=0
M1563 162 113 785 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=94450 $D=0
M1564 581 122 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=89820 $D=0
M1565 582 122 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=94450 $D=0
M1566 583 122 579 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=89820 $D=0
M1567 584 122 580 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=94450 $D=0
M1568 10 581 583 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=89820 $D=0
M1569 11 582 584 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=94450 $D=0
M1570 586 585 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=89820 $D=0
M1571 587 123 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=94450 $D=0
M1572 161 590 588 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=89820 $D=0
M1573 162 591 589 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=94450 $D=0
M1574 592 575 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=89820 $D=0
M1575 593 576 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=94450 $D=0
M1576 590 575 585 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=89820 $D=0
M1577 591 576 123 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=94450 $D=0
M1578 586 592 590 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=89820 $D=0
M1579 587 593 591 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=94450 $D=0
M1580 594 588 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=89820 $D=0
M1581 595 589 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=94450 $D=0
M1582 596 588 583 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=89820 $D=0
M1583 585 589 584 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=94450 $D=0
M1584 575 594 596 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=89820 $D=0
M1585 576 595 585 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=94450 $D=0
M1586 597 596 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=89820 $D=0
M1587 598 585 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=94450 $D=0
M1588 599 588 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=89820 $D=0
M1589 600 589 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=94450 $D=0
M1590 601 588 597 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=89820 $D=0
M1591 602 589 598 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=94450 $D=0
M1592 583 599 601 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=89820 $D=0
M1593 584 600 602 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=94450 $D=0
M1594 796 575 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=89460 $D=0
M1595 797 576 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=94090 $D=0
M1596 603 583 796 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=89460 $D=0
M1597 604 584 797 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=94090 $D=0
M1598 605 601 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=89820 $D=0
M1599 606 602 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=94450 $D=0
M1600 607 575 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=89820 $D=0
M1601 608 576 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=94450 $D=0
M1602 161 583 607 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=89820 $D=0
M1603 162 584 608 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=94450 $D=0
M1604 609 575 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=89820 $D=0
M1605 610 576 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=94450 $D=0
M1606 161 583 609 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=89820 $D=0
M1607 162 584 610 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=94450 $D=0
M1608 798 575 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=89640 $D=0
M1609 799 576 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=94270 $D=0
M1610 613 583 798 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=89640 $D=0
M1611 614 584 799 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=94270 $D=0
M1612 161 609 613 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=89820 $D=0
M1613 162 610 614 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=94450 $D=0
M1614 615 126 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=89820 $D=0
M1615 616 126 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=94450 $D=0
M1616 617 126 603 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=89820 $D=0
M1617 618 126 604 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=94450 $D=0
M1618 607 615 617 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=89820 $D=0
M1619 608 616 618 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=94450 $D=0
M1620 619 126 605 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=89820 $D=0
M1621 620 126 606 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=94450 $D=0
M1622 613 615 619 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=89820 $D=0
M1623 614 616 620 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=94450 $D=0
M1624 621 127 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=89820 $D=0
M1625 622 127 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=94450 $D=0
M1626 623 127 619 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=89820 $D=0
M1627 624 127 620 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=94450 $D=0
M1628 617 621 623 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=89820 $D=0
M1629 618 622 624 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=94450 $D=0
M1630 12 623 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=89820 $D=0
M1631 13 624 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=94450 $D=0
M1632 625 128 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=89820 $D=0
M1633 626 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=94450 $D=0
M1634 627 128 129 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=89820 $D=0
M1635 628 128 130 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=94450 $D=0
M1636 131 625 627 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=89820 $D=0
M1637 132 626 628 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=94450 $D=0
M1638 629 128 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=89820 $D=0
M1639 630 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=94450 $D=0
M1640 631 128 133 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=89820 $D=0
M1641 632 128 134 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=94450 $D=0
M1642 135 629 631 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=89820 $D=0
M1643 136 630 632 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=94450 $D=0
M1644 633 128 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=89820 $D=0
M1645 634 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=94450 $D=0
M1646 635 128 136 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=89820 $D=0
M1647 636 128 137 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=94450 $D=0
M1648 114 633 635 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=89820 $D=0
M1649 116 634 636 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=94450 $D=0
M1650 637 128 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=89820 $D=0
M1651 638 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=94450 $D=0
M1652 639 128 138 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=89820 $D=0
M1653 640 128 139 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=94450 $D=0
M1654 115 637 639 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=89820 $D=0
M1655 117 638 640 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=94450 $D=0
M1656 641 128 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=89820 $D=0
M1657 642 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=94450 $D=0
M1658 643 128 5 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=89820 $D=0
M1659 644 128 6 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=94450 $D=0
M1660 140 641 643 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=89820 $D=0
M1661 141 642 644 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=94450 $D=0
M1662 161 575 786 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=89820 $D=0
M1663 162 576 787 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=94450 $D=0
M1664 132 786 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=89820 $D=0
M1665 129 787 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=94450 $D=0
M1666 645 142 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=89820 $D=0
M1667 646 142 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=94450 $D=0
M1668 143 142 132 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=89820 $D=0
M1669 144 142 129 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=94450 $D=0
M1670 627 645 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=89820 $D=0
M1671 628 646 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=94450 $D=0
M1672 647 145 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=89820 $D=0
M1673 648 145 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=94450 $D=0
M1674 121 145 143 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=89820 $D=0
M1675 146 145 144 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=94450 $D=0
M1676 631 647 121 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=89820 $D=0
M1677 632 648 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=94450 $D=0
M1678 649 147 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=89820 $D=0
M1679 650 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=94450 $D=0
M1680 124 147 121 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=89820 $D=0
M1681 125 147 146 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=94450 $D=0
M1682 635 649 124 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=89820 $D=0
M1683 636 650 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=94450 $D=0
M1684 651 148 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=89820 $D=0
M1685 652 148 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=94450 $D=0
M1686 149 148 124 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=89820 $D=0
M1687 150 148 125 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=94450 $D=0
M1688 639 651 149 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=89820 $D=0
M1689 640 652 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=94450 $D=0
M1690 653 151 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=89820 $D=0
M1691 654 151 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=94450 $D=0
M1692 225 151 149 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=89820 $D=0
M1693 226 151 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=94450 $D=0
M1694 643 653 225 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=89820 $D=0
M1695 644 654 226 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=94450 $D=0
M1696 655 152 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=89820 $D=0
M1697 656 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=94450 $D=0
M1698 657 152 112 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=89820 $D=0
M1699 658 152 113 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=94450 $D=0
M1700 10 655 657 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=89820 $D=0
M1701 11 656 658 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=94450 $D=0
M1702 659 565 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=89820 $D=0
M1703 660 566 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=94450 $D=0
M1704 161 657 659 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=89820 $D=0
M1705 162 658 660 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=94450 $D=0
M1706 800 565 161 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=89640 $D=0
M1707 801 566 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=94270 $D=0
M1708 663 657 800 161 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=89640 $D=0
M1709 664 658 801 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=94270 $D=0
M1710 161 659 663 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=89820 $D=0
M1711 162 660 664 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=94450 $D=0
M1712 788 153 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=89820 $D=0
M1713 789 665 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=94450 $D=0
M1714 161 663 788 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=89820 $D=0
M1715 162 664 789 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=94450 $D=0
M1716 665 788 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=89820 $D=0
M1717 154 789 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=94450 $D=0
M1718 802 565 161 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=89460 $D=0
M1719 803 566 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=94090 $D=0
M1720 666 668 802 161 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=89460 $D=0
M1721 667 669 803 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=94090 $D=0
M1722 668 657 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=89820 $D=0
M1723 669 658 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=94450 $D=0
M1724 670 666 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=89820 $D=0
M1725 671 667 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=94450 $D=0
M1726 161 153 670 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=89820 $D=0
M1727 162 665 671 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=94450 $D=0
M1728 673 155 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=89820 $D=0
M1729 674 672 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=94450 $D=0
M1730 672 670 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=89820 $D=0
M1731 156 671 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=94450 $D=0
M1732 161 673 672 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=89820 $D=0
M1733 162 674 156 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=94450 $D=0
M1734 676 675 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=89820 $D=0
M1735 677 157 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=94450 $D=0
M1736 161 680 678 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=89820 $D=0
M1737 162 681 679 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=94450 $D=0
M1738 682 119 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=89820 $D=0
M1739 683 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=94450 $D=0
M1740 680 119 675 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=89820 $D=0
M1741 681 119 157 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=94450 $D=0
M1742 676 682 680 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=89820 $D=0
M1743 677 683 681 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=94450 $D=0
M1744 684 678 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=89820 $D=0
M1745 685 679 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=94450 $D=0
M1746 158 678 5 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=89820 $D=0
M1747 675 679 6 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=94450 $D=0
M1748 119 684 158 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=89820 $D=0
M1749 119 685 675 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=94450 $D=0
M1750 686 158 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=89820 $D=0
M1751 687 675 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=94450 $D=0
M1752 688 678 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=89820 $D=0
M1753 689 679 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=94450 $D=0
M1754 227 678 686 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=89820 $D=0
M1755 228 679 687 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=94450 $D=0
M1756 5 688 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=89820 $D=0
M1757 6 689 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=94450 $D=0
M1758 690 159 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=89820 $D=0
M1759 691 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=94450 $D=0
M1760 692 159 227 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=89820 $D=0
M1761 693 159 228 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=94450 $D=0
M1762 12 690 692 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=89820 $D=0
M1763 13 691 693 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=94450 $D=0
M1764 694 160 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=89820 $D=0
M1765 695 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=94450 $D=0
M1766 160 160 692 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=89820 $D=0
M1767 160 160 693 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=94450 $D=0
M1768 5 694 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=89820 $D=0
M1769 6 695 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=94450 $D=0
M1770 696 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=89820 $D=0
M1771 697 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=94450 $D=0
M1772 161 696 698 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=89820 $D=0
M1773 162 697 699 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=94450 $D=0
M1774 700 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=89820 $D=0
M1775 701 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=94450 $D=0
M1776 702 698 160 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=89820 $D=0
M1777 703 699 160 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=94450 $D=0
M1778 161 702 790 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=89820 $D=0
M1779 162 703 791 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=94450 $D=0
M1780 704 790 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=89820 $D=0
M1781 705 791 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=94450 $D=0
M1782 702 696 704 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=89820 $D=0
M1783 703 697 705 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=94450 $D=0
M1784 706 700 704 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=89820 $D=0
M1785 707 701 705 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=94450 $D=0
M1786 161 710 708 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=89820 $D=0
M1787 162 711 709 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=94450 $D=0
M1788 710 111 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=89820 $D=0
M1789 711 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=94450 $D=0
M1790 792 706 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=89820 $D=0
M1791 793 707 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=94450 $D=0
M1792 712 710 792 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=89820 $D=0
M1793 713 711 793 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=94450 $D=0
M1794 161 712 119 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=89820 $D=0
M1795 162 713 119 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=94450 $D=0
M1796 794 119 161 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=89820 $D=0
M1797 795 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=94450 $D=0
M1798 712 708 794 161 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=89820 $D=0
M1799 713 709 795 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=94450 $D=0
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163
** N=817 EP=163 IP=1514 FDC=1800
M0 203 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=79310 $D=1
M1 204 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=83940 $D=1
M2 205 203 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=79310 $D=1
M3 206 204 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=83940 $D=1
M4 5 1 205 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=79310 $D=1
M5 6 1 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=83940 $D=1
M6 207 203 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=79310 $D=1
M7 208 204 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=83940 $D=1
M8 2 1 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=79310 $D=1
M9 3 1 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=83940 $D=1
M10 209 203 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=79310 $D=1
M11 210 204 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=83940 $D=1
M12 2 1 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=79310 $D=1
M13 3 1 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=83940 $D=1
M14 213 211 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=79310 $D=1
M15 214 212 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=83940 $D=1
M16 211 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=79310 $D=1
M17 212 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=83940 $D=1
M18 215 211 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=79310 $D=1
M19 216 212 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=83940 $D=1
M20 205 7 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=79310 $D=1
M21 206 7 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=83940 $D=1
M22 217 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=79310 $D=1
M23 218 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=83940 $D=1
M24 219 217 215 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=79310 $D=1
M25 220 218 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=83940 $D=1
M26 213 8 219 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=79310 $D=1
M27 214 8 220 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=83940 $D=1
M28 221 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=79310 $D=1
M29 222 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=83940 $D=1
M30 223 221 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=79310 $D=1
M31 224 222 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=83940 $D=1
M32 10 9 223 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=79310 $D=1
M33 11 9 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=83940 $D=1
M34 225 221 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=79310 $D=1
M35 226 222 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=83940 $D=1
M36 227 9 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=79310 $D=1
M37 228 9 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=83940 $D=1
M38 231 221 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=79310 $D=1
M39 232 222 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=83940 $D=1
M40 219 9 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=79310 $D=1
M41 220 9 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=83940 $D=1
M42 235 233 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=79310 $D=1
M43 236 234 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=83940 $D=1
M44 233 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=79310 $D=1
M45 234 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=83940 $D=1
M46 237 233 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=79310 $D=1
M47 238 234 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=83940 $D=1
M48 223 14 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=79310 $D=1
M49 224 14 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=83940 $D=1
M50 239 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=79310 $D=1
M51 240 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=83940 $D=1
M52 241 239 237 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=79310 $D=1
M53 242 240 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=83940 $D=1
M54 235 15 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=79310 $D=1
M55 236 15 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=83940 $D=1
M56 5 16 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=79310 $D=1
M57 6 16 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=83940 $D=1
M58 245 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=79310 $D=1
M59 246 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=83940 $D=1
M60 247 16 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=79310 $D=1
M61 248 16 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=83940 $D=1
M62 5 247 716 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=79310 $D=1
M63 6 248 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=83940 $D=1
M64 249 716 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=79310 $D=1
M65 250 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=83940 $D=1
M66 247 243 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=79310 $D=1
M67 248 244 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=83940 $D=1
M68 249 17 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=79310 $D=1
M69 250 17 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=83940 $D=1
M70 255 18 249 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=79310 $D=1
M71 256 18 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=83940 $D=1
M72 253 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=79310 $D=1
M73 254 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=83940 $D=1
M74 5 19 257 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=79310 $D=1
M75 6 19 258 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=83940 $D=1
M76 259 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=79310 $D=1
M77 260 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=83940 $D=1
M78 261 19 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=79310 $D=1
M79 262 19 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=83940 $D=1
M80 5 261 718 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=79310 $D=1
M81 6 262 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=83940 $D=1
M82 263 718 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=79310 $D=1
M83 264 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=83940 $D=1
M84 261 257 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=79310 $D=1
M85 262 258 264 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=83940 $D=1
M86 263 20 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=79310 $D=1
M87 264 20 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=83940 $D=1
M88 255 21 263 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=79310 $D=1
M89 256 21 264 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=83940 $D=1
M90 265 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=79310 $D=1
M91 266 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=83940 $D=1
M92 5 22 267 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=79310 $D=1
M93 6 22 268 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=83940 $D=1
M94 269 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=79310 $D=1
M95 270 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=83940 $D=1
M96 271 22 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=79310 $D=1
M97 272 22 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=83940 $D=1
M98 5 271 720 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=79310 $D=1
M99 6 272 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=83940 $D=1
M100 273 720 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=79310 $D=1
M101 274 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=83940 $D=1
M102 271 267 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=79310 $D=1
M103 272 268 274 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=83940 $D=1
M104 273 23 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=79310 $D=1
M105 274 23 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=83940 $D=1
M106 255 24 273 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=79310 $D=1
M107 256 24 274 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=83940 $D=1
M108 275 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=79310 $D=1
M109 276 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=83940 $D=1
M110 5 25 277 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=79310 $D=1
M111 6 25 278 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=83940 $D=1
M112 279 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=79310 $D=1
M113 280 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=83940 $D=1
M114 281 25 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=79310 $D=1
M115 282 25 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=83940 $D=1
M116 5 281 722 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=79310 $D=1
M117 6 282 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=83940 $D=1
M118 283 722 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=79310 $D=1
M119 284 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=83940 $D=1
M120 281 277 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=79310 $D=1
M121 282 278 284 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=83940 $D=1
M122 283 26 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=79310 $D=1
M123 284 26 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=83940 $D=1
M124 255 27 283 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=79310 $D=1
M125 256 27 284 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=83940 $D=1
M126 285 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=79310 $D=1
M127 286 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=83940 $D=1
M128 5 28 287 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=79310 $D=1
M129 6 28 288 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=83940 $D=1
M130 289 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=79310 $D=1
M131 290 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=83940 $D=1
M132 291 28 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=79310 $D=1
M133 292 28 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=83940 $D=1
M134 5 291 724 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=79310 $D=1
M135 6 292 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=83940 $D=1
M136 293 724 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=79310 $D=1
M137 294 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=83940 $D=1
M138 291 287 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=79310 $D=1
M139 292 288 294 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=83940 $D=1
M140 293 29 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=79310 $D=1
M141 294 29 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=83940 $D=1
M142 255 30 293 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=79310 $D=1
M143 256 30 294 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=83940 $D=1
M144 295 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=79310 $D=1
M145 296 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=83940 $D=1
M146 5 31 297 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=79310 $D=1
M147 6 31 298 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=83940 $D=1
M148 299 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=79310 $D=1
M149 300 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=83940 $D=1
M150 301 31 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=79310 $D=1
M151 302 31 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=83940 $D=1
M152 5 301 726 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=79310 $D=1
M153 6 302 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=83940 $D=1
M154 303 726 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=79310 $D=1
M155 304 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=83940 $D=1
M156 301 297 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=79310 $D=1
M157 302 298 304 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=83940 $D=1
M158 303 32 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=79310 $D=1
M159 304 32 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=83940 $D=1
M160 255 33 303 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=79310 $D=1
M161 256 33 304 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=83940 $D=1
M162 305 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=79310 $D=1
M163 306 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=83940 $D=1
M164 5 34 307 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=79310 $D=1
M165 6 34 308 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=83940 $D=1
M166 309 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=79310 $D=1
M167 310 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=83940 $D=1
M168 311 34 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=79310 $D=1
M169 312 34 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=83940 $D=1
M170 5 311 728 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=79310 $D=1
M171 6 312 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=83940 $D=1
M172 313 728 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=79310 $D=1
M173 314 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=83940 $D=1
M174 311 307 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=79310 $D=1
M175 312 308 314 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=83940 $D=1
M176 313 35 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=79310 $D=1
M177 314 35 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=83940 $D=1
M178 255 36 313 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=79310 $D=1
M179 256 36 314 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=83940 $D=1
M180 315 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=79310 $D=1
M181 316 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=83940 $D=1
M182 5 37 317 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=79310 $D=1
M183 6 37 318 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=83940 $D=1
M184 319 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=79310 $D=1
M185 320 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=83940 $D=1
M186 321 37 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=79310 $D=1
M187 322 37 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=83940 $D=1
M188 5 321 730 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=79310 $D=1
M189 6 322 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=83940 $D=1
M190 323 730 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=79310 $D=1
M191 324 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=83940 $D=1
M192 321 317 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=79310 $D=1
M193 322 318 324 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=83940 $D=1
M194 323 38 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=79310 $D=1
M195 324 38 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=83940 $D=1
M196 255 39 323 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=79310 $D=1
M197 256 39 324 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=83940 $D=1
M198 325 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=79310 $D=1
M199 326 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=83940 $D=1
M200 5 40 327 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=79310 $D=1
M201 6 40 328 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=83940 $D=1
M202 329 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=79310 $D=1
M203 330 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=83940 $D=1
M204 331 40 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=79310 $D=1
M205 332 40 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=83940 $D=1
M206 5 331 732 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=79310 $D=1
M207 6 332 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=83940 $D=1
M208 333 732 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=79310 $D=1
M209 334 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=83940 $D=1
M210 331 327 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=79310 $D=1
M211 332 328 334 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=83940 $D=1
M212 333 41 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=79310 $D=1
M213 334 41 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=83940 $D=1
M214 255 42 333 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=79310 $D=1
M215 256 42 334 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=83940 $D=1
M216 335 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=79310 $D=1
M217 336 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=83940 $D=1
M218 5 43 337 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=79310 $D=1
M219 6 43 338 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=83940 $D=1
M220 339 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=79310 $D=1
M221 340 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=83940 $D=1
M222 341 43 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=79310 $D=1
M223 342 43 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=83940 $D=1
M224 5 341 734 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=79310 $D=1
M225 6 342 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=83940 $D=1
M226 343 734 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=79310 $D=1
M227 344 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=83940 $D=1
M228 341 337 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=79310 $D=1
M229 342 338 344 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=83940 $D=1
M230 343 44 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=79310 $D=1
M231 344 44 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=83940 $D=1
M232 255 45 343 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=79310 $D=1
M233 256 45 344 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=83940 $D=1
M234 345 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=79310 $D=1
M235 346 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=83940 $D=1
M236 5 46 347 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=79310 $D=1
M237 6 46 348 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=83940 $D=1
M238 349 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=79310 $D=1
M239 350 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=83940 $D=1
M240 351 46 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=79310 $D=1
M241 352 46 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=83940 $D=1
M242 5 351 736 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=79310 $D=1
M243 6 352 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=83940 $D=1
M244 353 736 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=79310 $D=1
M245 354 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=83940 $D=1
M246 351 347 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=79310 $D=1
M247 352 348 354 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=83940 $D=1
M248 353 47 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=79310 $D=1
M249 354 47 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=83940 $D=1
M250 255 48 353 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=79310 $D=1
M251 256 48 354 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=83940 $D=1
M252 355 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=79310 $D=1
M253 356 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=83940 $D=1
M254 5 49 357 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=79310 $D=1
M255 6 49 358 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=83940 $D=1
M256 359 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=79310 $D=1
M257 360 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=83940 $D=1
M258 361 49 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=79310 $D=1
M259 362 49 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=83940 $D=1
M260 5 361 738 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=79310 $D=1
M261 6 362 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=83940 $D=1
M262 363 738 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=79310 $D=1
M263 364 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=83940 $D=1
M264 361 357 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=79310 $D=1
M265 362 358 364 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=83940 $D=1
M266 363 50 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=79310 $D=1
M267 364 50 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=83940 $D=1
M268 255 51 363 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=79310 $D=1
M269 256 51 364 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=83940 $D=1
M270 365 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=79310 $D=1
M271 366 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=83940 $D=1
M272 5 52 367 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=79310 $D=1
M273 6 52 368 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=83940 $D=1
M274 369 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=79310 $D=1
M275 370 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=83940 $D=1
M276 371 52 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=79310 $D=1
M277 372 52 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=83940 $D=1
M278 5 371 740 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=79310 $D=1
M279 6 372 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=83940 $D=1
M280 373 740 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=79310 $D=1
M281 374 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=83940 $D=1
M282 371 367 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=79310 $D=1
M283 372 368 374 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=83940 $D=1
M284 373 53 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=79310 $D=1
M285 374 53 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=83940 $D=1
M286 255 54 373 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=79310 $D=1
M287 256 54 374 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=83940 $D=1
M288 375 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=79310 $D=1
M289 376 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=83940 $D=1
M290 5 55 377 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=79310 $D=1
M291 6 55 378 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=83940 $D=1
M292 379 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=79310 $D=1
M293 380 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=83940 $D=1
M294 381 55 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=79310 $D=1
M295 382 55 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=83940 $D=1
M296 5 381 742 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=79310 $D=1
M297 6 382 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=83940 $D=1
M298 383 742 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=79310 $D=1
M299 384 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=83940 $D=1
M300 381 377 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=79310 $D=1
M301 382 378 384 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=83940 $D=1
M302 383 56 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=79310 $D=1
M303 384 56 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=83940 $D=1
M304 255 57 383 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=79310 $D=1
M305 256 57 384 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=83940 $D=1
M306 385 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=79310 $D=1
M307 386 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=83940 $D=1
M308 5 58 387 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=79310 $D=1
M309 6 58 388 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=83940 $D=1
M310 389 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=79310 $D=1
M311 390 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=83940 $D=1
M312 391 58 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=79310 $D=1
M313 392 58 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=83940 $D=1
M314 5 391 744 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=79310 $D=1
M315 6 392 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=83940 $D=1
M316 393 744 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=79310 $D=1
M317 394 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=83940 $D=1
M318 391 387 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=79310 $D=1
M319 392 388 394 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=83940 $D=1
M320 393 59 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=79310 $D=1
M321 394 59 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=83940 $D=1
M322 255 60 393 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=79310 $D=1
M323 256 60 394 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=83940 $D=1
M324 395 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=79310 $D=1
M325 396 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=83940 $D=1
M326 5 61 397 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=79310 $D=1
M327 6 61 398 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=83940 $D=1
M328 399 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=79310 $D=1
M329 400 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=83940 $D=1
M330 401 61 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=79310 $D=1
M331 402 61 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=83940 $D=1
M332 5 401 746 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=79310 $D=1
M333 6 402 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=83940 $D=1
M334 403 746 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=79310 $D=1
M335 404 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=83940 $D=1
M336 401 397 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=79310 $D=1
M337 402 398 404 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=83940 $D=1
M338 403 62 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=79310 $D=1
M339 404 62 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=83940 $D=1
M340 255 63 403 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=79310 $D=1
M341 256 63 404 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=83940 $D=1
M342 405 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=79310 $D=1
M343 406 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=83940 $D=1
M344 5 64 407 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=79310 $D=1
M345 6 64 408 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=83940 $D=1
M346 409 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=79310 $D=1
M347 410 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=83940 $D=1
M348 411 64 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=79310 $D=1
M349 412 64 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=83940 $D=1
M350 5 411 748 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=79310 $D=1
M351 6 412 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=83940 $D=1
M352 413 748 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=79310 $D=1
M353 414 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=83940 $D=1
M354 411 407 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=79310 $D=1
M355 412 408 414 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=83940 $D=1
M356 413 65 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=79310 $D=1
M357 414 65 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=83940 $D=1
M358 255 66 413 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=79310 $D=1
M359 256 66 414 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=83940 $D=1
M360 415 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=79310 $D=1
M361 416 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=83940 $D=1
M362 5 67 417 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=79310 $D=1
M363 6 67 418 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=83940 $D=1
M364 419 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=79310 $D=1
M365 420 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=83940 $D=1
M366 421 67 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=79310 $D=1
M367 422 67 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=83940 $D=1
M368 5 421 750 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=79310 $D=1
M369 6 422 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=83940 $D=1
M370 423 750 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=79310 $D=1
M371 424 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=83940 $D=1
M372 421 417 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=79310 $D=1
M373 422 418 424 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=83940 $D=1
M374 423 68 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=79310 $D=1
M375 424 68 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=83940 $D=1
M376 255 69 423 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=79310 $D=1
M377 256 69 424 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=83940 $D=1
M378 425 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=79310 $D=1
M379 426 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=83940 $D=1
M380 5 70 427 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=79310 $D=1
M381 6 70 428 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=83940 $D=1
M382 429 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=79310 $D=1
M383 430 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=83940 $D=1
M384 431 70 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=79310 $D=1
M385 432 70 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=83940 $D=1
M386 5 431 752 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=79310 $D=1
M387 6 432 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=83940 $D=1
M388 433 752 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=79310 $D=1
M389 434 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=83940 $D=1
M390 431 427 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=79310 $D=1
M391 432 428 434 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=83940 $D=1
M392 433 71 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=79310 $D=1
M393 434 71 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=83940 $D=1
M394 255 72 433 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=79310 $D=1
M395 256 72 434 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=83940 $D=1
M396 435 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=79310 $D=1
M397 436 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=83940 $D=1
M398 5 73 437 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=79310 $D=1
M399 6 73 438 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=83940 $D=1
M400 439 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=79310 $D=1
M401 440 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=83940 $D=1
M402 441 73 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=79310 $D=1
M403 442 73 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=83940 $D=1
M404 5 441 754 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=79310 $D=1
M405 6 442 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=83940 $D=1
M406 443 754 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=79310 $D=1
M407 444 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=83940 $D=1
M408 441 437 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=79310 $D=1
M409 442 438 444 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=83940 $D=1
M410 443 74 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=79310 $D=1
M411 444 74 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=83940 $D=1
M412 255 75 443 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=79310 $D=1
M413 256 75 444 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=83940 $D=1
M414 445 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=79310 $D=1
M415 446 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=83940 $D=1
M416 5 76 447 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=79310 $D=1
M417 6 76 448 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=83940 $D=1
M418 449 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=79310 $D=1
M419 450 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=83940 $D=1
M420 451 76 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=79310 $D=1
M421 452 76 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=83940 $D=1
M422 5 451 756 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=79310 $D=1
M423 6 452 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=83940 $D=1
M424 453 756 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=79310 $D=1
M425 454 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=83940 $D=1
M426 451 447 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=79310 $D=1
M427 452 448 454 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=83940 $D=1
M428 453 77 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=79310 $D=1
M429 454 77 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=83940 $D=1
M430 255 78 453 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=79310 $D=1
M431 256 78 454 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=83940 $D=1
M432 455 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=79310 $D=1
M433 456 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=83940 $D=1
M434 5 79 457 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=79310 $D=1
M435 6 79 458 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=83940 $D=1
M436 459 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=79310 $D=1
M437 460 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=83940 $D=1
M438 461 79 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=79310 $D=1
M439 462 79 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=83940 $D=1
M440 5 461 758 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=79310 $D=1
M441 6 462 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=83940 $D=1
M442 463 758 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=79310 $D=1
M443 464 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=83940 $D=1
M444 461 457 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=79310 $D=1
M445 462 458 464 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=83940 $D=1
M446 463 80 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=79310 $D=1
M447 464 80 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=83940 $D=1
M448 255 81 463 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=79310 $D=1
M449 256 81 464 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=83940 $D=1
M450 465 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=79310 $D=1
M451 466 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=83940 $D=1
M452 5 82 467 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=79310 $D=1
M453 6 82 468 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=83940 $D=1
M454 469 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=79310 $D=1
M455 470 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=83940 $D=1
M456 471 82 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=79310 $D=1
M457 472 82 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=83940 $D=1
M458 5 471 760 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=79310 $D=1
M459 6 472 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=83940 $D=1
M460 473 760 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=79310 $D=1
M461 474 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=83940 $D=1
M462 471 467 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=79310 $D=1
M463 472 468 474 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=83940 $D=1
M464 473 83 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=79310 $D=1
M465 474 83 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=83940 $D=1
M466 255 84 473 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=79310 $D=1
M467 256 84 474 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=83940 $D=1
M468 475 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=79310 $D=1
M469 476 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=83940 $D=1
M470 5 85 477 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=79310 $D=1
M471 6 85 478 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=83940 $D=1
M472 479 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=79310 $D=1
M473 480 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=83940 $D=1
M474 481 85 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=79310 $D=1
M475 482 85 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=83940 $D=1
M476 5 481 762 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=79310 $D=1
M477 6 482 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=83940 $D=1
M478 483 762 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=79310 $D=1
M479 484 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=83940 $D=1
M480 481 477 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=79310 $D=1
M481 482 478 484 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=83940 $D=1
M482 483 86 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=79310 $D=1
M483 484 86 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=83940 $D=1
M484 255 87 483 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=79310 $D=1
M485 256 87 484 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=83940 $D=1
M486 485 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=79310 $D=1
M487 486 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=83940 $D=1
M488 5 88 487 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=79310 $D=1
M489 6 88 488 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=83940 $D=1
M490 489 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=79310 $D=1
M491 490 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=83940 $D=1
M492 491 88 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=79310 $D=1
M493 492 88 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=83940 $D=1
M494 5 491 764 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=79310 $D=1
M495 6 492 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=83940 $D=1
M496 493 764 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=79310 $D=1
M497 494 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=83940 $D=1
M498 491 487 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=79310 $D=1
M499 492 488 494 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=83940 $D=1
M500 493 89 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=79310 $D=1
M501 494 89 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=83940 $D=1
M502 255 90 493 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=79310 $D=1
M503 256 90 494 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=83940 $D=1
M504 495 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=79310 $D=1
M505 496 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=83940 $D=1
M506 5 91 497 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=79310 $D=1
M507 6 91 498 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=83940 $D=1
M508 499 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=79310 $D=1
M509 500 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=83940 $D=1
M510 501 91 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=79310 $D=1
M511 502 91 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=83940 $D=1
M512 5 501 766 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=79310 $D=1
M513 6 502 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=83940 $D=1
M514 503 766 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=79310 $D=1
M515 504 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=83940 $D=1
M516 501 497 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=79310 $D=1
M517 502 498 504 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=83940 $D=1
M518 503 92 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=79310 $D=1
M519 504 92 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=83940 $D=1
M520 255 93 503 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=79310 $D=1
M521 256 93 504 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=83940 $D=1
M522 505 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=79310 $D=1
M523 506 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=83940 $D=1
M524 5 94 507 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=79310 $D=1
M525 6 94 508 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=83940 $D=1
M526 509 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=79310 $D=1
M527 510 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=83940 $D=1
M528 511 94 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=79310 $D=1
M529 512 94 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=83940 $D=1
M530 5 511 768 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=79310 $D=1
M531 6 512 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=83940 $D=1
M532 513 768 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=79310 $D=1
M533 514 769 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=83940 $D=1
M534 511 507 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=79310 $D=1
M535 512 508 514 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=83940 $D=1
M536 513 95 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=79310 $D=1
M537 514 95 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=83940 $D=1
M538 255 96 513 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=79310 $D=1
M539 256 96 514 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=83940 $D=1
M540 515 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=79310 $D=1
M541 516 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=83940 $D=1
M542 5 97 517 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=79310 $D=1
M543 6 97 518 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=83940 $D=1
M544 519 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=79310 $D=1
M545 520 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=83940 $D=1
M546 521 97 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=79310 $D=1
M547 522 97 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=83940 $D=1
M548 5 521 770 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=79310 $D=1
M549 6 522 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=83940 $D=1
M550 523 770 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=79310 $D=1
M551 524 771 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=83940 $D=1
M552 521 517 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=79310 $D=1
M553 522 518 524 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=83940 $D=1
M554 523 98 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=79310 $D=1
M555 524 98 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=83940 $D=1
M556 255 99 523 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=79310 $D=1
M557 256 99 524 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=83940 $D=1
M558 525 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=79310 $D=1
M559 526 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=83940 $D=1
M560 5 100 527 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=79310 $D=1
M561 6 100 528 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=83940 $D=1
M562 529 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=79310 $D=1
M563 530 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=83940 $D=1
M564 531 100 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=79310 $D=1
M565 532 100 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=83940 $D=1
M566 5 531 772 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=79310 $D=1
M567 6 532 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=83940 $D=1
M568 533 772 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=79310 $D=1
M569 534 773 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=83940 $D=1
M570 531 527 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=79310 $D=1
M571 532 528 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=83940 $D=1
M572 533 101 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=79310 $D=1
M573 534 101 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=83940 $D=1
M574 255 102 533 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=79310 $D=1
M575 256 102 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=83940 $D=1
M576 535 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=79310 $D=1
M577 536 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=83940 $D=1
M578 5 103 537 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=79310 $D=1
M579 6 103 538 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=83940 $D=1
M580 539 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=79310 $D=1
M581 540 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=83940 $D=1
M582 541 103 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=79310 $D=1
M583 542 103 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=83940 $D=1
M584 5 541 774 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=79310 $D=1
M585 6 542 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=83940 $D=1
M586 543 774 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=79310 $D=1
M587 544 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=83940 $D=1
M588 541 537 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=79310 $D=1
M589 542 538 544 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=83940 $D=1
M590 543 104 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=79310 $D=1
M591 544 104 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=83940 $D=1
M592 255 105 543 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=79310 $D=1
M593 256 105 544 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=83940 $D=1
M594 545 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=79310 $D=1
M595 546 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=83940 $D=1
M596 5 106 547 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=79310 $D=1
M597 6 106 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=83940 $D=1
M598 549 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=79310 $D=1
M599 550 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=83940 $D=1
M600 551 106 241 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=79310 $D=1
M601 552 106 242 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=83940 $D=1
M602 5 551 776 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=79310 $D=1
M603 6 552 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=83940 $D=1
M604 553 776 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=79310 $D=1
M605 554 777 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=83940 $D=1
M606 551 547 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=79310 $D=1
M607 552 548 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=83940 $D=1
M608 553 107 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=79310 $D=1
M609 554 107 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=83940 $D=1
M610 255 108 553 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=79310 $D=1
M611 256 108 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=83940 $D=1
M612 555 108 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=79310 $D=1
M613 556 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=83940 $D=1
M614 5 109 557 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=79310 $D=1
M615 6 109 558 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=83940 $D=1
M616 559 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=79310 $D=1
M617 560 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=83940 $D=1
M618 5 110 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=79310 $D=1
M619 6 110 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=83940 $D=1
M620 255 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=79310 $D=1
M621 256 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=83940 $D=1
M622 5 563 561 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=79310 $D=1
M623 6 564 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=83940 $D=1
M624 563 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=79310 $D=1
M625 564 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=83940 $D=1
M626 778 251 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=79310 $D=1
M627 779 252 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=83940 $D=1
M628 565 561 778 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=79310 $D=1
M629 566 562 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=83940 $D=1
M630 5 565 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=79310 $D=1
M631 6 566 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=83940 $D=1
M632 780 567 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=79310 $D=1
M633 781 568 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=83940 $D=1
M634 565 563 780 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=79310 $D=1
M635 566 564 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=83940 $D=1
M636 5 572 570 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=79310 $D=1
M637 6 573 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=83940 $D=1
M638 572 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=79310 $D=1
M639 573 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=83940 $D=1
M640 782 255 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=79310 $D=1
M641 783 256 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=83940 $D=1
M642 574 570 782 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=79310 $D=1
M643 575 571 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=83940 $D=1
M644 5 574 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=79310 $D=1
M645 6 575 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=83940 $D=1
M646 784 117 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=79310 $D=1
M647 785 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=83940 $D=1
M648 574 572 784 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=79310 $D=1
M649 575 573 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=83940 $D=1
M650 576 119 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=79310 $D=1
M651 577 119 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=83940 $D=1
M652 578 576 567 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=79310 $D=1
M653 579 577 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=83940 $D=1
M654 121 119 578 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=79310 $D=1
M655 121 119 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=83940 $D=1
M656 580 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=79310 $D=1
M657 581 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=83940 $D=1
M658 582 580 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=79310 $D=1
M659 583 581 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=83940 $D=1
M660 786 122 582 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=79310 $D=1
M661 787 122 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=83940 $D=1
M662 5 117 786 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=79310 $D=1
M663 6 118 787 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=83940 $D=1
M664 584 124 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=79310 $D=1
M665 585 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=83940 $D=1
M666 586 584 582 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=79310 $D=1
M667 587 585 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=83940 $D=1
M668 10 124 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=79310 $D=1
M669 11 124 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=83940 $D=1
M670 589 588 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=79310 $D=1
M671 590 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=83940 $D=1
M672 5 593 591 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=79310 $D=1
M673 6 594 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=83940 $D=1
M674 595 578 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=79310 $D=1
M675 596 579 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=83940 $D=1
M676 593 595 588 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=79310 $D=1
M677 594 596 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=83940 $D=1
M678 589 578 593 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=79310 $D=1
M679 590 579 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=83940 $D=1
M680 597 591 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=79310 $D=1
M681 598 592 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=83940 $D=1
M682 127 597 586 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=79310 $D=1
M683 588 598 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=83940 $D=1
M684 578 591 127 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=79310 $D=1
M685 579 592 588 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=83940 $D=1
M686 599 127 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=79310 $D=1
M687 600 588 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=83940 $D=1
M688 601 591 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=79310 $D=1
M689 602 592 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=83940 $D=1
M690 603 601 599 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=79310 $D=1
M691 604 602 600 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=83940 $D=1
M692 586 591 603 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=79310 $D=1
M693 587 592 604 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=83940 $D=1
M694 605 578 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=79310 $D=1
M695 606 579 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=83940 $D=1
M696 5 586 605 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=79310 $D=1
M697 6 587 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=83940 $D=1
M698 607 603 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=79310 $D=1
M699 608 604 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=83940 $D=1
M700 806 578 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=79310 $D=1
M701 807 579 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=83940 $D=1
M702 609 586 806 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=79310 $D=1
M703 610 587 807 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=83940 $D=1
M704 808 578 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=79310 $D=1
M705 809 579 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=83940 $D=1
M706 611 586 808 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=79310 $D=1
M707 612 587 809 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=83940 $D=1
M708 615 578 613 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=79310 $D=1
M709 616 579 614 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=83940 $D=1
M710 613 586 615 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=79310 $D=1
M711 614 587 616 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=83940 $D=1
M712 5 611 613 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=79310 $D=1
M713 6 612 614 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=83940 $D=1
M714 617 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=79310 $D=1
M715 618 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=83940 $D=1
M716 619 617 605 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=79310 $D=1
M717 620 618 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=83940 $D=1
M718 609 128 619 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=79310 $D=1
M719 610 128 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=83940 $D=1
M720 621 617 607 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=79310 $D=1
M721 622 618 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=83940 $D=1
M722 615 128 621 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=79310 $D=1
M723 616 128 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=83940 $D=1
M724 623 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=79310 $D=1
M725 624 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=83940 $D=1
M726 625 623 621 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=79310 $D=1
M727 626 624 622 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=83940 $D=1
M728 619 129 625 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=79310 $D=1
M729 620 129 626 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=83940 $D=1
M730 12 625 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=79310 $D=1
M731 13 626 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=83940 $D=1
M732 627 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=79310 $D=1
M733 628 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=83940 $D=1
M734 629 627 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=79310 $D=1
M735 630 628 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=83940 $D=1
M736 133 130 629 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=79310 $D=1
M737 134 130 630 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=83940 $D=1
M738 631 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=79310 $D=1
M739 632 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=83940 $D=1
M740 633 631 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=79310 $D=1
M741 634 632 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=83940 $D=1
M742 137 130 633 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=79310 $D=1
M743 138 130 634 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=83940 $D=1
M744 635 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=79310 $D=1
M745 636 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=83940 $D=1
M746 637 635 138 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=79310 $D=1
M747 638 636 139 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=83940 $D=1
M748 113 130 637 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=79310 $D=1
M749 115 130 638 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=83940 $D=1
M750 639 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=79310 $D=1
M751 640 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=83940 $D=1
M752 641 639 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=79310 $D=1
M753 642 640 141 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=83940 $D=1
M754 114 130 641 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=79310 $D=1
M755 116 130 642 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=83940 $D=1
M756 643 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=79310 $D=1
M757 644 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=83940 $D=1
M758 645 643 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=79310 $D=1
M759 646 644 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=83940 $D=1
M760 142 130 645 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=79310 $D=1
M761 143 130 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=83940 $D=1
M762 5 578 788 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=79310 $D=1
M763 6 579 789 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=83940 $D=1
M764 134 788 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=79310 $D=1
M765 131 789 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=83940 $D=1
M766 647 144 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=79310 $D=1
M767 648 144 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=83940 $D=1
M768 145 647 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=79310 $D=1
M769 146 648 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=83940 $D=1
M770 629 144 145 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=79310 $D=1
M771 630 144 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=83940 $D=1
M772 649 147 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=79310 $D=1
M773 650 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=83940 $D=1
M774 120 649 145 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=79310 $D=1
M775 123 650 146 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=83940 $D=1
M776 633 147 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=79310 $D=1
M777 634 147 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=83940 $D=1
M778 651 148 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=79310 $D=1
M779 652 148 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=83940 $D=1
M780 112 651 120 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=79310 $D=1
M781 126 652 123 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=83940 $D=1
M782 637 148 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=79310 $D=1
M783 638 148 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=83940 $D=1
M784 653 149 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=79310 $D=1
M785 654 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=83940 $D=1
M786 150 653 112 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=79310 $D=1
M787 151 654 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=83940 $D=1
M788 641 149 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=79310 $D=1
M789 642 149 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=83940 $D=1
M790 655 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=79310 $D=1
M791 656 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=83940 $D=1
M792 227 655 150 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=79310 $D=1
M793 228 656 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=83940 $D=1
M794 645 152 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=79310 $D=1
M795 646 152 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=83940 $D=1
M796 657 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=79310 $D=1
M797 658 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=83940 $D=1
M798 659 657 117 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=79310 $D=1
M799 660 658 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=83940 $D=1
M800 10 153 659 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=79310 $D=1
M801 11 153 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=83940 $D=1
M802 810 567 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=79310 $D=1
M803 811 568 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=83940 $D=1
M804 661 659 810 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=79310 $D=1
M805 662 660 811 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=83940 $D=1
M806 665 567 663 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=79310 $D=1
M807 666 568 664 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=83940 $D=1
M808 663 659 665 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=79310 $D=1
M809 664 660 666 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=83940 $D=1
M810 5 661 663 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=79310 $D=1
M811 6 662 664 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=83940 $D=1
M812 812 154 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=79310 $D=1
M813 813 667 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=83940 $D=1
M814 790 665 812 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=79310 $D=1
M815 791 666 813 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=83940 $D=1
M816 667 790 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=79310 $D=1
M817 155 791 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=83940 $D=1
M818 668 567 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=79310 $D=1
M819 669 568 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=83940 $D=1
M820 5 670 668 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=79310 $D=1
M821 6 671 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=83940 $D=1
M822 670 659 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=79310 $D=1
M823 671 660 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=83940 $D=1
M824 814 668 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=79310 $D=1
M825 815 669 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=83940 $D=1
M826 672 154 814 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=79310 $D=1
M827 673 667 815 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=83940 $D=1
M828 675 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=79310 $D=1
M829 676 674 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=83940 $D=1
M830 816 672 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=79310 $D=1
M831 817 673 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=83940 $D=1
M832 674 675 816 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=79310 $D=1
M833 157 676 817 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=83940 $D=1
M834 678 677 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=79310 $D=1
M835 679 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=83940 $D=1
M836 5 682 680 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=79310 $D=1
M837 6 683 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=83940 $D=1
M838 684 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=79310 $D=1
M839 685 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=83940 $D=1
M840 682 684 677 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=79310 $D=1
M841 683 685 158 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=83940 $D=1
M842 678 121 682 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=79310 $D=1
M843 679 121 683 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=83940 $D=1
M844 686 680 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=79310 $D=1
M845 687 681 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=83940 $D=1
M846 159 686 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=79310 $D=1
M847 677 687 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=83940 $D=1
M848 121 680 159 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=79310 $D=1
M849 121 681 677 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=83940 $D=1
M850 688 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=79310 $D=1
M851 689 677 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=83940 $D=1
M852 690 680 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=79310 $D=1
M853 691 681 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=83940 $D=1
M854 229 690 688 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=79310 $D=1
M855 230 691 689 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=83940 $D=1
M856 5 680 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=79310 $D=1
M857 6 681 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=83940 $D=1
M858 692 160 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=79310 $D=1
M859 693 160 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=83940 $D=1
M860 694 692 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=79310 $D=1
M861 695 693 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=83940 $D=1
M862 12 160 694 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=79310 $D=1
M863 13 160 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=83940 $D=1
M864 696 161 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=79310 $D=1
M865 697 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=83940 $D=1
M866 161 696 694 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=79310 $D=1
M867 161 697 695 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=83940 $D=1
M868 5 161 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=79310 $D=1
M869 6 161 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=83940 $D=1
M870 698 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=79310 $D=1
M871 699 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=83940 $D=1
M872 5 698 700 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=79310 $D=1
M873 6 699 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=83940 $D=1
M874 702 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=79310 $D=1
M875 703 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=83940 $D=1
M876 704 698 161 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=79310 $D=1
M877 705 699 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=83940 $D=1
M878 5 704 792 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=79310 $D=1
M879 6 705 793 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=83940 $D=1
M880 706 792 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=79310 $D=1
M881 707 793 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=83940 $D=1
M882 704 700 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=79310 $D=1
M883 705 701 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=83940 $D=1
M884 708 111 706 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=79310 $D=1
M885 709 111 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=83940 $D=1
M886 5 712 710 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=79310 $D=1
M887 6 713 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=83940 $D=1
M888 712 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=79310 $D=1
M889 713 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=83940 $D=1
M890 794 708 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=79310 $D=1
M891 795 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=83940 $D=1
M892 714 710 794 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=79310 $D=1
M893 715 711 795 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=83940 $D=1
M894 5 714 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=79310 $D=1
M895 6 715 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=83940 $D=1
M896 796 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=79310 $D=1
M897 797 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=83940 $D=1
M898 714 712 796 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=79310 $D=1
M899 715 713 797 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=83940 $D=1
M900 203 1 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=80560 $D=0
M901 204 1 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=85190 $D=0
M902 205 1 2 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=80560 $D=0
M903 206 1 3 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=85190 $D=0
M904 5 203 205 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=80560 $D=0
M905 6 204 206 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=85190 $D=0
M906 207 1 4 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=80560 $D=0
M907 208 1 4 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=85190 $D=0
M908 2 203 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=80560 $D=0
M909 3 204 208 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=85190 $D=0
M910 209 1 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=80560 $D=0
M911 210 1 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=85190 $D=0
M912 2 203 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=80560 $D=0
M913 3 204 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=85190 $D=0
M914 213 7 209 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=80560 $D=0
M915 214 7 210 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=85190 $D=0
M916 211 7 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=80560 $D=0
M917 212 7 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=85190 $D=0
M918 215 7 207 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=80560 $D=0
M919 216 7 208 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=85190 $D=0
M920 205 211 215 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=80560 $D=0
M921 206 212 216 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=85190 $D=0
M922 217 8 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=80560 $D=0
M923 218 8 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=85190 $D=0
M924 219 8 215 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=80560 $D=0
M925 220 8 216 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=85190 $D=0
M926 213 217 219 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=80560 $D=0
M927 214 218 220 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=85190 $D=0
M928 221 9 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=80560 $D=0
M929 222 9 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=85190 $D=0
M930 223 9 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=80560 $D=0
M931 224 9 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=85190 $D=0
M932 10 221 223 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=80560 $D=0
M933 11 222 224 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=85190 $D=0
M934 225 9 12 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=80560 $D=0
M935 226 9 13 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=85190 $D=0
M936 227 221 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=80560 $D=0
M937 228 222 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=85190 $D=0
M938 231 9 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=80560 $D=0
M939 232 9 230 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=85190 $D=0
M940 219 221 231 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=80560 $D=0
M941 220 222 232 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=85190 $D=0
M942 235 14 231 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=80560 $D=0
M943 236 14 232 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=85190 $D=0
M944 233 14 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=80560 $D=0
M945 234 14 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=85190 $D=0
M946 237 14 225 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=80560 $D=0
M947 238 14 226 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=85190 $D=0
M948 223 233 237 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=80560 $D=0
M949 224 234 238 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=85190 $D=0
M950 239 15 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=80560 $D=0
M951 240 15 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=85190 $D=0
M952 241 15 237 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=80560 $D=0
M953 242 15 238 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=85190 $D=0
M954 235 239 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=80560 $D=0
M955 236 240 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=85190 $D=0
M956 162 16 243 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=80560 $D=0
M957 163 16 244 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=85190 $D=0
M958 245 17 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=80560 $D=0
M959 246 17 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=85190 $D=0
M960 247 243 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=80560 $D=0
M961 248 244 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=85190 $D=0
M962 162 247 716 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=80560 $D=0
M963 163 248 717 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=85190 $D=0
M964 249 716 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=80560 $D=0
M965 250 717 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=85190 $D=0
M966 247 16 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=80560 $D=0
M967 248 16 250 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=85190 $D=0
M968 249 245 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=80560 $D=0
M969 250 246 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=85190 $D=0
M970 255 253 249 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=80560 $D=0
M971 256 254 250 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=85190 $D=0
M972 253 18 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=80560 $D=0
M973 254 18 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=85190 $D=0
M974 162 19 257 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=80560 $D=0
M975 163 19 258 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=85190 $D=0
M976 259 20 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=80560 $D=0
M977 260 20 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=85190 $D=0
M978 261 257 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=80560 $D=0
M979 262 258 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=85190 $D=0
M980 162 261 718 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=80560 $D=0
M981 163 262 719 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=85190 $D=0
M982 263 718 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=80560 $D=0
M983 264 719 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=85190 $D=0
M984 261 19 263 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=80560 $D=0
M985 262 19 264 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=85190 $D=0
M986 263 259 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=80560 $D=0
M987 264 260 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=85190 $D=0
M988 255 265 263 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=80560 $D=0
M989 256 266 264 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=85190 $D=0
M990 265 21 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=80560 $D=0
M991 266 21 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=85190 $D=0
M992 162 22 267 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=80560 $D=0
M993 163 22 268 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=85190 $D=0
M994 269 23 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=80560 $D=0
M995 270 23 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=85190 $D=0
M996 271 267 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=80560 $D=0
M997 272 268 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=85190 $D=0
M998 162 271 720 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=80560 $D=0
M999 163 272 721 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=85190 $D=0
M1000 273 720 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=80560 $D=0
M1001 274 721 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=85190 $D=0
M1002 271 22 273 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=80560 $D=0
M1003 272 22 274 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=85190 $D=0
M1004 273 269 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=80560 $D=0
M1005 274 270 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=85190 $D=0
M1006 255 275 273 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=80560 $D=0
M1007 256 276 274 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=85190 $D=0
M1008 275 24 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=80560 $D=0
M1009 276 24 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=85190 $D=0
M1010 162 25 277 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=80560 $D=0
M1011 163 25 278 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=85190 $D=0
M1012 279 26 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=80560 $D=0
M1013 280 26 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=85190 $D=0
M1014 281 277 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=80560 $D=0
M1015 282 278 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=85190 $D=0
M1016 162 281 722 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=80560 $D=0
M1017 163 282 723 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=85190 $D=0
M1018 283 722 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=80560 $D=0
M1019 284 723 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=85190 $D=0
M1020 281 25 283 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=80560 $D=0
M1021 282 25 284 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=85190 $D=0
M1022 283 279 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=80560 $D=0
M1023 284 280 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=85190 $D=0
M1024 255 285 283 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=80560 $D=0
M1025 256 286 284 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=85190 $D=0
M1026 285 27 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=80560 $D=0
M1027 286 27 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=85190 $D=0
M1028 162 28 287 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=80560 $D=0
M1029 163 28 288 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=85190 $D=0
M1030 289 29 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=80560 $D=0
M1031 290 29 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=85190 $D=0
M1032 291 287 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=80560 $D=0
M1033 292 288 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=85190 $D=0
M1034 162 291 724 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=80560 $D=0
M1035 163 292 725 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=85190 $D=0
M1036 293 724 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=80560 $D=0
M1037 294 725 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=85190 $D=0
M1038 291 28 293 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=80560 $D=0
M1039 292 28 294 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=85190 $D=0
M1040 293 289 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=80560 $D=0
M1041 294 290 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=85190 $D=0
M1042 255 295 293 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=80560 $D=0
M1043 256 296 294 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=85190 $D=0
M1044 295 30 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=80560 $D=0
M1045 296 30 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=85190 $D=0
M1046 162 31 297 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=80560 $D=0
M1047 163 31 298 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=85190 $D=0
M1048 299 32 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=80560 $D=0
M1049 300 32 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=85190 $D=0
M1050 301 297 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=80560 $D=0
M1051 302 298 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=85190 $D=0
M1052 162 301 726 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=80560 $D=0
M1053 163 302 727 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=85190 $D=0
M1054 303 726 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=80560 $D=0
M1055 304 727 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=85190 $D=0
M1056 301 31 303 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=80560 $D=0
M1057 302 31 304 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=85190 $D=0
M1058 303 299 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=80560 $D=0
M1059 304 300 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=85190 $D=0
M1060 255 305 303 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=80560 $D=0
M1061 256 306 304 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=85190 $D=0
M1062 305 33 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=80560 $D=0
M1063 306 33 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=85190 $D=0
M1064 162 34 307 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=80560 $D=0
M1065 163 34 308 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=85190 $D=0
M1066 309 35 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=80560 $D=0
M1067 310 35 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=85190 $D=0
M1068 311 307 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=80560 $D=0
M1069 312 308 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=85190 $D=0
M1070 162 311 728 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=80560 $D=0
M1071 163 312 729 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=85190 $D=0
M1072 313 728 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=80560 $D=0
M1073 314 729 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=85190 $D=0
M1074 311 34 313 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=80560 $D=0
M1075 312 34 314 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=85190 $D=0
M1076 313 309 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=80560 $D=0
M1077 314 310 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=85190 $D=0
M1078 255 315 313 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=80560 $D=0
M1079 256 316 314 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=85190 $D=0
M1080 315 36 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=80560 $D=0
M1081 316 36 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=85190 $D=0
M1082 162 37 317 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=80560 $D=0
M1083 163 37 318 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=85190 $D=0
M1084 319 38 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=80560 $D=0
M1085 320 38 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=85190 $D=0
M1086 321 317 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=80560 $D=0
M1087 322 318 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=85190 $D=0
M1088 162 321 730 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=80560 $D=0
M1089 163 322 731 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=85190 $D=0
M1090 323 730 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=80560 $D=0
M1091 324 731 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=85190 $D=0
M1092 321 37 323 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=80560 $D=0
M1093 322 37 324 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=85190 $D=0
M1094 323 319 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=80560 $D=0
M1095 324 320 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=85190 $D=0
M1096 255 325 323 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=80560 $D=0
M1097 256 326 324 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=85190 $D=0
M1098 325 39 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=80560 $D=0
M1099 326 39 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=85190 $D=0
M1100 162 40 327 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=80560 $D=0
M1101 163 40 328 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=85190 $D=0
M1102 329 41 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=80560 $D=0
M1103 330 41 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=85190 $D=0
M1104 331 327 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=80560 $D=0
M1105 332 328 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=85190 $D=0
M1106 162 331 732 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=80560 $D=0
M1107 163 332 733 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=85190 $D=0
M1108 333 732 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=80560 $D=0
M1109 334 733 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=85190 $D=0
M1110 331 40 333 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=80560 $D=0
M1111 332 40 334 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=85190 $D=0
M1112 333 329 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=80560 $D=0
M1113 334 330 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=85190 $D=0
M1114 255 335 333 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=80560 $D=0
M1115 256 336 334 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=85190 $D=0
M1116 335 42 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=80560 $D=0
M1117 336 42 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=85190 $D=0
M1118 162 43 337 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=80560 $D=0
M1119 163 43 338 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=85190 $D=0
M1120 339 44 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=80560 $D=0
M1121 340 44 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=85190 $D=0
M1122 341 337 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=80560 $D=0
M1123 342 338 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=85190 $D=0
M1124 162 341 734 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=80560 $D=0
M1125 163 342 735 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=85190 $D=0
M1126 343 734 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=80560 $D=0
M1127 344 735 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=85190 $D=0
M1128 341 43 343 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=80560 $D=0
M1129 342 43 344 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=85190 $D=0
M1130 343 339 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=80560 $D=0
M1131 344 340 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=85190 $D=0
M1132 255 345 343 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=80560 $D=0
M1133 256 346 344 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=85190 $D=0
M1134 345 45 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=80560 $D=0
M1135 346 45 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=85190 $D=0
M1136 162 46 347 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=80560 $D=0
M1137 163 46 348 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=85190 $D=0
M1138 349 47 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=80560 $D=0
M1139 350 47 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=85190 $D=0
M1140 351 347 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=80560 $D=0
M1141 352 348 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=85190 $D=0
M1142 162 351 736 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=80560 $D=0
M1143 163 352 737 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=85190 $D=0
M1144 353 736 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=80560 $D=0
M1145 354 737 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=85190 $D=0
M1146 351 46 353 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=80560 $D=0
M1147 352 46 354 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=85190 $D=0
M1148 353 349 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=80560 $D=0
M1149 354 350 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=85190 $D=0
M1150 255 355 353 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=80560 $D=0
M1151 256 356 354 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=85190 $D=0
M1152 355 48 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=80560 $D=0
M1153 356 48 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=85190 $D=0
M1154 162 49 357 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=80560 $D=0
M1155 163 49 358 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=85190 $D=0
M1156 359 50 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=80560 $D=0
M1157 360 50 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=85190 $D=0
M1158 361 357 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=80560 $D=0
M1159 362 358 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=85190 $D=0
M1160 162 361 738 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=80560 $D=0
M1161 163 362 739 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=85190 $D=0
M1162 363 738 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=80560 $D=0
M1163 364 739 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=85190 $D=0
M1164 361 49 363 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=80560 $D=0
M1165 362 49 364 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=85190 $D=0
M1166 363 359 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=80560 $D=0
M1167 364 360 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=85190 $D=0
M1168 255 365 363 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=80560 $D=0
M1169 256 366 364 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=85190 $D=0
M1170 365 51 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=80560 $D=0
M1171 366 51 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=85190 $D=0
M1172 162 52 367 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=80560 $D=0
M1173 163 52 368 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=85190 $D=0
M1174 369 53 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=80560 $D=0
M1175 370 53 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=85190 $D=0
M1176 371 367 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=80560 $D=0
M1177 372 368 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=85190 $D=0
M1178 162 371 740 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=80560 $D=0
M1179 163 372 741 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=85190 $D=0
M1180 373 740 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=80560 $D=0
M1181 374 741 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=85190 $D=0
M1182 371 52 373 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=80560 $D=0
M1183 372 52 374 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=85190 $D=0
M1184 373 369 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=80560 $D=0
M1185 374 370 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=85190 $D=0
M1186 255 375 373 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=80560 $D=0
M1187 256 376 374 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=85190 $D=0
M1188 375 54 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=80560 $D=0
M1189 376 54 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=85190 $D=0
M1190 162 55 377 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=80560 $D=0
M1191 163 55 378 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=85190 $D=0
M1192 379 56 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=80560 $D=0
M1193 380 56 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=85190 $D=0
M1194 381 377 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=80560 $D=0
M1195 382 378 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=85190 $D=0
M1196 162 381 742 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=80560 $D=0
M1197 163 382 743 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=85190 $D=0
M1198 383 742 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=80560 $D=0
M1199 384 743 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=85190 $D=0
M1200 381 55 383 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=80560 $D=0
M1201 382 55 384 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=85190 $D=0
M1202 383 379 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=80560 $D=0
M1203 384 380 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=85190 $D=0
M1204 255 385 383 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=80560 $D=0
M1205 256 386 384 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=85190 $D=0
M1206 385 57 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=80560 $D=0
M1207 386 57 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=85190 $D=0
M1208 162 58 387 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=80560 $D=0
M1209 163 58 388 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=85190 $D=0
M1210 389 59 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=80560 $D=0
M1211 390 59 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=85190 $D=0
M1212 391 387 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=80560 $D=0
M1213 392 388 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=85190 $D=0
M1214 162 391 744 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=80560 $D=0
M1215 163 392 745 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=85190 $D=0
M1216 393 744 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=80560 $D=0
M1217 394 745 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=85190 $D=0
M1218 391 58 393 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=80560 $D=0
M1219 392 58 394 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=85190 $D=0
M1220 393 389 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=80560 $D=0
M1221 394 390 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=85190 $D=0
M1222 255 395 393 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=80560 $D=0
M1223 256 396 394 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=85190 $D=0
M1224 395 60 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=80560 $D=0
M1225 396 60 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=85190 $D=0
M1226 162 61 397 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=80560 $D=0
M1227 163 61 398 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=85190 $D=0
M1228 399 62 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=80560 $D=0
M1229 400 62 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=85190 $D=0
M1230 401 397 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=80560 $D=0
M1231 402 398 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=85190 $D=0
M1232 162 401 746 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=80560 $D=0
M1233 163 402 747 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=85190 $D=0
M1234 403 746 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=80560 $D=0
M1235 404 747 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=85190 $D=0
M1236 401 61 403 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=80560 $D=0
M1237 402 61 404 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=85190 $D=0
M1238 403 399 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=80560 $D=0
M1239 404 400 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=85190 $D=0
M1240 255 405 403 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=80560 $D=0
M1241 256 406 404 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=85190 $D=0
M1242 405 63 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=80560 $D=0
M1243 406 63 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=85190 $D=0
M1244 162 64 407 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=80560 $D=0
M1245 163 64 408 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=85190 $D=0
M1246 409 65 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=80560 $D=0
M1247 410 65 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=85190 $D=0
M1248 411 407 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=80560 $D=0
M1249 412 408 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=85190 $D=0
M1250 162 411 748 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=80560 $D=0
M1251 163 412 749 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=85190 $D=0
M1252 413 748 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=80560 $D=0
M1253 414 749 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=85190 $D=0
M1254 411 64 413 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=80560 $D=0
M1255 412 64 414 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=85190 $D=0
M1256 413 409 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=80560 $D=0
M1257 414 410 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=85190 $D=0
M1258 255 415 413 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=80560 $D=0
M1259 256 416 414 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=85190 $D=0
M1260 415 66 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=80560 $D=0
M1261 416 66 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=85190 $D=0
M1262 162 67 417 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=80560 $D=0
M1263 163 67 418 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=85190 $D=0
M1264 419 68 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=80560 $D=0
M1265 420 68 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=85190 $D=0
M1266 421 417 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=80560 $D=0
M1267 422 418 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=85190 $D=0
M1268 162 421 750 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=80560 $D=0
M1269 163 422 751 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=85190 $D=0
M1270 423 750 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=80560 $D=0
M1271 424 751 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=85190 $D=0
M1272 421 67 423 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=80560 $D=0
M1273 422 67 424 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=85190 $D=0
M1274 423 419 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=80560 $D=0
M1275 424 420 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=85190 $D=0
M1276 255 425 423 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=80560 $D=0
M1277 256 426 424 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=85190 $D=0
M1278 425 69 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=80560 $D=0
M1279 426 69 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=85190 $D=0
M1280 162 70 427 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=80560 $D=0
M1281 163 70 428 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=85190 $D=0
M1282 429 71 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=80560 $D=0
M1283 430 71 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=85190 $D=0
M1284 431 427 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=80560 $D=0
M1285 432 428 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=85190 $D=0
M1286 162 431 752 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=80560 $D=0
M1287 163 432 753 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=85190 $D=0
M1288 433 752 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=80560 $D=0
M1289 434 753 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=85190 $D=0
M1290 431 70 433 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=80560 $D=0
M1291 432 70 434 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=85190 $D=0
M1292 433 429 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=80560 $D=0
M1293 434 430 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=85190 $D=0
M1294 255 435 433 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=80560 $D=0
M1295 256 436 434 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=85190 $D=0
M1296 435 72 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=80560 $D=0
M1297 436 72 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=85190 $D=0
M1298 162 73 437 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=80560 $D=0
M1299 163 73 438 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=85190 $D=0
M1300 439 74 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=80560 $D=0
M1301 440 74 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=85190 $D=0
M1302 441 437 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=80560 $D=0
M1303 442 438 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=85190 $D=0
M1304 162 441 754 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=80560 $D=0
M1305 163 442 755 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=85190 $D=0
M1306 443 754 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=80560 $D=0
M1307 444 755 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=85190 $D=0
M1308 441 73 443 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=80560 $D=0
M1309 442 73 444 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=85190 $D=0
M1310 443 439 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=80560 $D=0
M1311 444 440 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=85190 $D=0
M1312 255 445 443 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=80560 $D=0
M1313 256 446 444 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=85190 $D=0
M1314 445 75 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=80560 $D=0
M1315 446 75 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=85190 $D=0
M1316 162 76 447 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=80560 $D=0
M1317 163 76 448 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=85190 $D=0
M1318 449 77 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=80560 $D=0
M1319 450 77 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=85190 $D=0
M1320 451 447 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=80560 $D=0
M1321 452 448 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=85190 $D=0
M1322 162 451 756 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=80560 $D=0
M1323 163 452 757 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=85190 $D=0
M1324 453 756 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=80560 $D=0
M1325 454 757 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=85190 $D=0
M1326 451 76 453 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=80560 $D=0
M1327 452 76 454 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=85190 $D=0
M1328 453 449 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=80560 $D=0
M1329 454 450 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=85190 $D=0
M1330 255 455 453 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=80560 $D=0
M1331 256 456 454 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=85190 $D=0
M1332 455 78 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=80560 $D=0
M1333 456 78 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=85190 $D=0
M1334 162 79 457 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=80560 $D=0
M1335 163 79 458 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=85190 $D=0
M1336 459 80 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=80560 $D=0
M1337 460 80 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=85190 $D=0
M1338 461 457 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=80560 $D=0
M1339 462 458 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=85190 $D=0
M1340 162 461 758 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=80560 $D=0
M1341 163 462 759 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=85190 $D=0
M1342 463 758 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=80560 $D=0
M1343 464 759 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=85190 $D=0
M1344 461 79 463 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=80560 $D=0
M1345 462 79 464 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=85190 $D=0
M1346 463 459 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=80560 $D=0
M1347 464 460 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=85190 $D=0
M1348 255 465 463 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=80560 $D=0
M1349 256 466 464 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=85190 $D=0
M1350 465 81 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=80560 $D=0
M1351 466 81 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=85190 $D=0
M1352 162 82 467 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=80560 $D=0
M1353 163 82 468 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=85190 $D=0
M1354 469 83 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=80560 $D=0
M1355 470 83 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=85190 $D=0
M1356 471 467 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=80560 $D=0
M1357 472 468 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=85190 $D=0
M1358 162 471 760 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=80560 $D=0
M1359 163 472 761 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=85190 $D=0
M1360 473 760 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=80560 $D=0
M1361 474 761 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=85190 $D=0
M1362 471 82 473 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=80560 $D=0
M1363 472 82 474 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=85190 $D=0
M1364 473 469 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=80560 $D=0
M1365 474 470 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=85190 $D=0
M1366 255 475 473 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=80560 $D=0
M1367 256 476 474 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=85190 $D=0
M1368 475 84 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=80560 $D=0
M1369 476 84 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=85190 $D=0
M1370 162 85 477 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=80560 $D=0
M1371 163 85 478 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=85190 $D=0
M1372 479 86 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=80560 $D=0
M1373 480 86 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=85190 $D=0
M1374 481 477 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=80560 $D=0
M1375 482 478 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=85190 $D=0
M1376 162 481 762 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=80560 $D=0
M1377 163 482 763 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=85190 $D=0
M1378 483 762 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=80560 $D=0
M1379 484 763 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=85190 $D=0
M1380 481 85 483 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=80560 $D=0
M1381 482 85 484 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=85190 $D=0
M1382 483 479 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=80560 $D=0
M1383 484 480 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=85190 $D=0
M1384 255 485 483 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=80560 $D=0
M1385 256 486 484 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=85190 $D=0
M1386 485 87 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=80560 $D=0
M1387 486 87 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=85190 $D=0
M1388 162 88 487 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=80560 $D=0
M1389 163 88 488 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=85190 $D=0
M1390 489 89 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=80560 $D=0
M1391 490 89 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=85190 $D=0
M1392 491 487 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=80560 $D=0
M1393 492 488 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=85190 $D=0
M1394 162 491 764 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=80560 $D=0
M1395 163 492 765 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=85190 $D=0
M1396 493 764 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=80560 $D=0
M1397 494 765 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=85190 $D=0
M1398 491 88 493 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=80560 $D=0
M1399 492 88 494 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=85190 $D=0
M1400 493 489 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=80560 $D=0
M1401 494 490 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=85190 $D=0
M1402 255 495 493 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=80560 $D=0
M1403 256 496 494 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=85190 $D=0
M1404 495 90 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=80560 $D=0
M1405 496 90 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=85190 $D=0
M1406 162 91 497 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=80560 $D=0
M1407 163 91 498 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=85190 $D=0
M1408 499 92 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=80560 $D=0
M1409 500 92 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=85190 $D=0
M1410 501 497 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=80560 $D=0
M1411 502 498 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=85190 $D=0
M1412 162 501 766 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=80560 $D=0
M1413 163 502 767 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=85190 $D=0
M1414 503 766 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=80560 $D=0
M1415 504 767 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=85190 $D=0
M1416 501 91 503 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=80560 $D=0
M1417 502 91 504 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=85190 $D=0
M1418 503 499 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=80560 $D=0
M1419 504 500 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=85190 $D=0
M1420 255 505 503 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=80560 $D=0
M1421 256 506 504 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=85190 $D=0
M1422 505 93 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=80560 $D=0
M1423 506 93 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=85190 $D=0
M1424 162 94 507 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=80560 $D=0
M1425 163 94 508 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=85190 $D=0
M1426 509 95 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=80560 $D=0
M1427 510 95 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=85190 $D=0
M1428 511 507 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=80560 $D=0
M1429 512 508 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=85190 $D=0
M1430 162 511 768 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=80560 $D=0
M1431 163 512 769 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=85190 $D=0
M1432 513 768 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=80560 $D=0
M1433 514 769 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=85190 $D=0
M1434 511 94 513 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=80560 $D=0
M1435 512 94 514 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=85190 $D=0
M1436 513 509 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=80560 $D=0
M1437 514 510 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=85190 $D=0
M1438 255 515 513 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=80560 $D=0
M1439 256 516 514 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=85190 $D=0
M1440 515 96 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=80560 $D=0
M1441 516 96 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=85190 $D=0
M1442 162 97 517 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=80560 $D=0
M1443 163 97 518 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=85190 $D=0
M1444 519 98 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=80560 $D=0
M1445 520 98 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=85190 $D=0
M1446 521 517 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=80560 $D=0
M1447 522 518 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=85190 $D=0
M1448 162 521 770 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=80560 $D=0
M1449 163 522 771 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=85190 $D=0
M1450 523 770 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=80560 $D=0
M1451 524 771 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=85190 $D=0
M1452 521 97 523 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=80560 $D=0
M1453 522 97 524 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=85190 $D=0
M1454 523 519 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=80560 $D=0
M1455 524 520 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=85190 $D=0
M1456 255 525 523 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=80560 $D=0
M1457 256 526 524 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=85190 $D=0
M1458 525 99 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=80560 $D=0
M1459 526 99 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=85190 $D=0
M1460 162 100 527 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=80560 $D=0
M1461 163 100 528 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=85190 $D=0
M1462 529 101 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=80560 $D=0
M1463 530 101 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=85190 $D=0
M1464 531 527 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=80560 $D=0
M1465 532 528 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=85190 $D=0
M1466 162 531 772 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=80560 $D=0
M1467 163 532 773 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=85190 $D=0
M1468 533 772 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=80560 $D=0
M1469 534 773 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=85190 $D=0
M1470 531 100 533 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=80560 $D=0
M1471 532 100 534 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=85190 $D=0
M1472 533 529 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=80560 $D=0
M1473 534 530 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=85190 $D=0
M1474 255 535 533 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=80560 $D=0
M1475 256 536 534 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=85190 $D=0
M1476 535 102 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=80560 $D=0
M1477 536 102 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=85190 $D=0
M1478 162 103 537 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=80560 $D=0
M1479 163 103 538 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=85190 $D=0
M1480 539 104 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=80560 $D=0
M1481 540 104 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=85190 $D=0
M1482 541 537 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=80560 $D=0
M1483 542 538 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=85190 $D=0
M1484 162 541 774 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=80560 $D=0
M1485 163 542 775 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=85190 $D=0
M1486 543 774 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=80560 $D=0
M1487 544 775 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=85190 $D=0
M1488 541 103 543 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=80560 $D=0
M1489 542 103 544 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=85190 $D=0
M1490 543 539 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=80560 $D=0
M1491 544 540 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=85190 $D=0
M1492 255 545 543 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=80560 $D=0
M1493 256 546 544 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=85190 $D=0
M1494 545 105 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=80560 $D=0
M1495 546 105 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=85190 $D=0
M1496 162 106 547 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=80560 $D=0
M1497 163 106 548 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=85190 $D=0
M1498 549 107 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=80560 $D=0
M1499 550 107 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=85190 $D=0
M1500 551 547 241 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=80560 $D=0
M1501 552 548 242 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=85190 $D=0
M1502 162 551 776 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=80560 $D=0
M1503 163 552 777 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=85190 $D=0
M1504 553 776 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=80560 $D=0
M1505 554 777 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=85190 $D=0
M1506 551 106 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=80560 $D=0
M1507 552 106 554 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=85190 $D=0
M1508 553 549 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=80560 $D=0
M1509 554 550 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=85190 $D=0
M1510 255 555 553 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=80560 $D=0
M1511 256 556 554 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=85190 $D=0
M1512 555 108 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=80560 $D=0
M1513 556 108 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=85190 $D=0
M1514 162 109 557 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=80560 $D=0
M1515 163 109 558 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=85190 $D=0
M1516 559 110 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=80560 $D=0
M1517 560 110 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=85190 $D=0
M1518 5 559 251 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=80560 $D=0
M1519 6 560 252 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=85190 $D=0
M1520 255 557 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=80560 $D=0
M1521 256 558 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=85190 $D=0
M1522 162 563 561 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=80560 $D=0
M1523 163 564 562 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=85190 $D=0
M1524 563 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=80560 $D=0
M1525 564 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=85190 $D=0
M1526 778 251 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=80560 $D=0
M1527 779 252 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=85190 $D=0
M1528 565 563 778 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=80560 $D=0
M1529 566 564 779 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=85190 $D=0
M1530 162 565 567 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=80560 $D=0
M1531 163 566 568 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=85190 $D=0
M1532 780 567 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=80560 $D=0
M1533 781 568 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=85190 $D=0
M1534 565 561 780 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=80560 $D=0
M1535 566 562 781 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=85190 $D=0
M1536 162 572 570 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=80560 $D=0
M1537 163 573 571 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=85190 $D=0
M1538 572 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=80560 $D=0
M1539 573 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=85190 $D=0
M1540 782 255 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=80560 $D=0
M1541 783 256 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=85190 $D=0
M1542 574 572 782 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=80560 $D=0
M1543 575 573 783 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=85190 $D=0
M1544 162 574 117 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=80560 $D=0
M1545 163 575 118 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=85190 $D=0
M1546 784 117 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=80560 $D=0
M1547 785 118 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=85190 $D=0
M1548 574 570 784 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=80560 $D=0
M1549 575 571 785 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=85190 $D=0
M1550 576 119 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=80560 $D=0
M1551 577 119 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=85190 $D=0
M1552 578 119 567 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=80560 $D=0
M1553 579 119 568 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=85190 $D=0
M1554 121 576 578 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=80560 $D=0
M1555 121 577 579 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=85190 $D=0
M1556 580 122 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=80560 $D=0
M1557 581 122 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=85190 $D=0
M1558 582 122 117 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=80560 $D=0
M1559 583 122 118 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=85190 $D=0
M1560 786 580 582 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=80560 $D=0
M1561 787 581 583 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=85190 $D=0
M1562 162 117 786 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=80560 $D=0
M1563 163 118 787 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=85190 $D=0
M1564 584 124 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=80560 $D=0
M1565 585 124 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=85190 $D=0
M1566 586 124 582 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=80560 $D=0
M1567 587 124 583 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=85190 $D=0
M1568 10 584 586 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=80560 $D=0
M1569 11 585 587 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=85190 $D=0
M1570 589 588 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=80560 $D=0
M1571 590 125 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=85190 $D=0
M1572 162 593 591 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=80560 $D=0
M1573 163 594 592 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=85190 $D=0
M1574 595 578 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=80560 $D=0
M1575 596 579 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=85190 $D=0
M1576 593 578 588 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=80560 $D=0
M1577 594 579 125 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=85190 $D=0
M1578 589 595 593 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=80560 $D=0
M1579 590 596 594 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=85190 $D=0
M1580 597 591 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=80560 $D=0
M1581 598 592 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=85190 $D=0
M1582 127 591 586 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=80560 $D=0
M1583 588 592 587 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=85190 $D=0
M1584 578 597 127 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=80560 $D=0
M1585 579 598 588 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=85190 $D=0
M1586 599 127 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=80560 $D=0
M1587 600 588 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=85190 $D=0
M1588 601 591 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=80560 $D=0
M1589 602 592 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=85190 $D=0
M1590 603 591 599 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=80560 $D=0
M1591 604 592 600 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=85190 $D=0
M1592 586 601 603 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=80560 $D=0
M1593 587 602 604 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=85190 $D=0
M1594 798 578 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=80200 $D=0
M1595 799 579 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=84830 $D=0
M1596 605 586 798 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=80200 $D=0
M1597 606 587 799 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=84830 $D=0
M1598 607 603 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=80560 $D=0
M1599 608 604 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=85190 $D=0
M1600 609 578 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=80560 $D=0
M1601 610 579 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=85190 $D=0
M1602 162 586 609 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=80560 $D=0
M1603 163 587 610 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=85190 $D=0
M1604 611 578 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=80560 $D=0
M1605 612 579 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=85190 $D=0
M1606 162 586 611 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=80560 $D=0
M1607 163 587 612 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=85190 $D=0
M1608 800 578 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=80380 $D=0
M1609 801 579 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=85010 $D=0
M1610 615 586 800 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=80380 $D=0
M1611 616 587 801 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=85010 $D=0
M1612 162 611 615 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=80560 $D=0
M1613 163 612 616 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=85190 $D=0
M1614 617 128 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=80560 $D=0
M1615 618 128 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=85190 $D=0
M1616 619 128 605 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=80560 $D=0
M1617 620 128 606 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=85190 $D=0
M1618 609 617 619 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=80560 $D=0
M1619 610 618 620 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=85190 $D=0
M1620 621 128 607 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=80560 $D=0
M1621 622 128 608 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=85190 $D=0
M1622 615 617 621 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=80560 $D=0
M1623 616 618 622 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=85190 $D=0
M1624 623 129 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=80560 $D=0
M1625 624 129 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=85190 $D=0
M1626 625 129 621 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=80560 $D=0
M1627 626 129 622 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=85190 $D=0
M1628 619 623 625 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=80560 $D=0
M1629 620 624 626 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=85190 $D=0
M1630 12 625 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=80560 $D=0
M1631 13 626 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=85190 $D=0
M1632 627 130 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=80560 $D=0
M1633 628 130 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=85190 $D=0
M1634 629 130 131 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=80560 $D=0
M1635 630 130 132 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=85190 $D=0
M1636 133 627 629 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=80560 $D=0
M1637 134 628 630 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=85190 $D=0
M1638 631 130 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=80560 $D=0
M1639 632 130 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=85190 $D=0
M1640 633 130 135 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=80560 $D=0
M1641 634 130 136 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=85190 $D=0
M1642 137 631 633 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=80560 $D=0
M1643 138 632 634 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=85190 $D=0
M1644 635 130 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=80560 $D=0
M1645 636 130 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=85190 $D=0
M1646 637 130 138 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=80560 $D=0
M1647 638 130 139 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=85190 $D=0
M1648 113 635 637 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=80560 $D=0
M1649 115 636 638 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=85190 $D=0
M1650 639 130 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=80560 $D=0
M1651 640 130 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=85190 $D=0
M1652 641 130 140 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=80560 $D=0
M1653 642 130 141 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=85190 $D=0
M1654 114 639 641 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=80560 $D=0
M1655 116 640 642 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=85190 $D=0
M1656 643 130 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=80560 $D=0
M1657 644 130 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=85190 $D=0
M1658 645 130 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=80560 $D=0
M1659 646 130 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=85190 $D=0
M1660 142 643 645 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=80560 $D=0
M1661 143 644 646 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=85190 $D=0
M1662 162 578 788 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=80560 $D=0
M1663 163 579 789 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=85190 $D=0
M1664 134 788 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=80560 $D=0
M1665 131 789 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=85190 $D=0
M1666 647 144 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=80560 $D=0
M1667 648 144 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=85190 $D=0
M1668 145 144 134 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=80560 $D=0
M1669 146 144 131 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=85190 $D=0
M1670 629 647 145 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=80560 $D=0
M1671 630 648 146 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=85190 $D=0
M1672 649 147 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=80560 $D=0
M1673 650 147 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=85190 $D=0
M1674 120 147 145 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=80560 $D=0
M1675 123 147 146 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=85190 $D=0
M1676 633 649 120 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=80560 $D=0
M1677 634 650 123 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=85190 $D=0
M1678 651 148 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=80560 $D=0
M1679 652 148 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=85190 $D=0
M1680 112 148 120 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=80560 $D=0
M1681 126 148 123 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=85190 $D=0
M1682 637 651 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=80560 $D=0
M1683 638 652 126 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=85190 $D=0
M1684 653 149 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=80560 $D=0
M1685 654 149 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=85190 $D=0
M1686 150 149 112 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=80560 $D=0
M1687 151 149 126 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=85190 $D=0
M1688 641 653 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=80560 $D=0
M1689 642 654 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=85190 $D=0
M1690 655 152 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=80560 $D=0
M1691 656 152 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=85190 $D=0
M1692 227 152 150 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=80560 $D=0
M1693 228 152 151 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=85190 $D=0
M1694 645 655 227 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=80560 $D=0
M1695 646 656 228 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=85190 $D=0
M1696 657 153 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=80560 $D=0
M1697 658 153 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=85190 $D=0
M1698 659 153 117 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=80560 $D=0
M1699 660 153 118 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=85190 $D=0
M1700 10 657 659 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=80560 $D=0
M1701 11 658 660 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=85190 $D=0
M1702 661 567 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=80560 $D=0
M1703 662 568 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=85190 $D=0
M1704 162 659 661 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=80560 $D=0
M1705 163 660 662 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=85190 $D=0
M1706 802 567 162 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=80380 $D=0
M1707 803 568 163 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=85010 $D=0
M1708 665 659 802 162 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=80380 $D=0
M1709 666 660 803 163 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=85010 $D=0
M1710 162 661 665 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=80560 $D=0
M1711 163 662 666 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=85190 $D=0
M1712 790 154 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=80560 $D=0
M1713 791 667 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=85190 $D=0
M1714 162 665 790 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=80560 $D=0
M1715 163 666 791 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=85190 $D=0
M1716 667 790 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=80560 $D=0
M1717 155 791 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=85190 $D=0
M1718 804 567 162 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=80200 $D=0
M1719 805 568 163 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=84830 $D=0
M1720 668 670 804 162 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=80200 $D=0
M1721 669 671 805 163 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=84830 $D=0
M1722 670 659 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=80560 $D=0
M1723 671 660 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=85190 $D=0
M1724 672 668 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=80560 $D=0
M1725 673 669 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=85190 $D=0
M1726 162 154 672 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=80560 $D=0
M1727 163 667 673 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=85190 $D=0
M1728 675 156 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=80560 $D=0
M1729 676 674 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=85190 $D=0
M1730 674 672 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=80560 $D=0
M1731 157 673 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=85190 $D=0
M1732 162 675 674 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=80560 $D=0
M1733 163 676 157 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=85190 $D=0
M1734 678 677 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=80560 $D=0
M1735 679 158 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=85190 $D=0
M1736 162 682 680 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=80560 $D=0
M1737 163 683 681 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=85190 $D=0
M1738 684 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=80560 $D=0
M1739 685 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=85190 $D=0
M1740 682 121 677 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=80560 $D=0
M1741 683 121 158 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=85190 $D=0
M1742 678 684 682 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=80560 $D=0
M1743 679 685 683 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=85190 $D=0
M1744 686 680 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=80560 $D=0
M1745 687 681 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=85190 $D=0
M1746 159 680 5 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=80560 $D=0
M1747 677 681 6 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=85190 $D=0
M1748 121 686 159 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=80560 $D=0
M1749 121 687 677 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=85190 $D=0
M1750 688 159 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=80560 $D=0
M1751 689 677 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=85190 $D=0
M1752 690 680 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=80560 $D=0
M1753 691 681 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=85190 $D=0
M1754 229 680 688 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=80560 $D=0
M1755 230 681 689 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=85190 $D=0
M1756 5 690 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=80560 $D=0
M1757 6 691 230 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=85190 $D=0
M1758 692 160 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=80560 $D=0
M1759 693 160 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=85190 $D=0
M1760 694 160 229 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=80560 $D=0
M1761 695 160 230 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=85190 $D=0
M1762 12 692 694 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=80560 $D=0
M1763 13 693 695 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=85190 $D=0
M1764 696 161 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=80560 $D=0
M1765 697 161 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=85190 $D=0
M1766 161 161 694 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=80560 $D=0
M1767 161 161 695 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=85190 $D=0
M1768 5 696 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=80560 $D=0
M1769 6 697 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=85190 $D=0
M1770 698 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=80560 $D=0
M1771 699 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=85190 $D=0
M1772 162 698 700 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=80560 $D=0
M1773 163 699 701 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=85190 $D=0
M1774 702 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=80560 $D=0
M1775 703 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=85190 $D=0
M1776 704 700 161 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=80560 $D=0
M1777 705 701 161 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=85190 $D=0
M1778 162 704 792 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=80560 $D=0
M1779 163 705 793 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=85190 $D=0
M1780 706 792 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=80560 $D=0
M1781 707 793 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=85190 $D=0
M1782 704 698 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=80560 $D=0
M1783 705 699 707 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=85190 $D=0
M1784 708 702 706 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=80560 $D=0
M1785 709 703 707 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=85190 $D=0
M1786 162 712 710 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=80560 $D=0
M1787 163 713 711 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=85190 $D=0
M1788 712 111 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=80560 $D=0
M1789 713 111 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=85190 $D=0
M1790 794 708 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=80560 $D=0
M1791 795 709 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=85190 $D=0
M1792 714 712 794 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=80560 $D=0
M1793 715 713 795 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=85190 $D=0
M1794 162 714 121 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=80560 $D=0
M1795 163 715 121 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=85190 $D=0
M1796 796 121 162 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=80560 $D=0
M1797 797 121 163 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=85190 $D=0
M1798 714 710 796 162 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=80560 $D=0
M1799 715 711 797 163 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=85190 $D=0
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166
** N=818 EP=165 IP=1514 FDC=1800
M0 205 1 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=70050 $D=1
M1 206 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=74680 $D=1
M2 207 205 2 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=70050 $D=1
M3 208 206 3 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=74680 $D=1
M4 5 1 207 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=70050 $D=1
M5 6 1 208 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=74680 $D=1
M6 209 205 4 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=70050 $D=1
M7 210 206 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=74680 $D=1
M8 3 1 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=70050 $D=1
M9 3 1 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=74680 $D=1
M10 211 205 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=70050 $D=1
M11 212 206 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=74680 $D=1
M12 5 1 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=70050 $D=1
M13 3 1 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=74680 $D=1
M14 215 213 211 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=70050 $D=1
M15 216 214 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=74680 $D=1
M16 213 7 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=70050 $D=1
M17 214 7 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=74680 $D=1
M18 217 213 209 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=70050 $D=1
M19 218 214 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=74680 $D=1
M20 207 7 217 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=70050 $D=1
M21 208 7 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=74680 $D=1
M22 219 8 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=70050 $D=1
M23 220 8 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=74680 $D=1
M24 221 219 217 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=70050 $D=1
M25 222 220 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=74680 $D=1
M26 215 8 221 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=70050 $D=1
M27 216 8 222 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=74680 $D=1
M28 223 9 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=70050 $D=1
M29 224 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=74680 $D=1
M30 225 223 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=70050 $D=1
M31 226 224 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=74680 $D=1
M32 10 9 225 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=70050 $D=1
M33 11 9 226 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=74680 $D=1
M34 227 223 12 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=70050 $D=1
M35 228 224 13 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=74680 $D=1
M36 229 9 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=70050 $D=1
M37 230 9 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=74680 $D=1
M38 233 223 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=70050 $D=1
M39 234 224 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=74680 $D=1
M40 221 9 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=70050 $D=1
M41 222 9 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=74680 $D=1
M42 237 235 233 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=70050 $D=1
M43 238 236 234 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=74680 $D=1
M44 235 14 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=70050 $D=1
M45 236 14 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=74680 $D=1
M46 239 235 227 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=70050 $D=1
M47 240 236 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=74680 $D=1
M48 225 14 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=70050 $D=1
M49 226 14 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=74680 $D=1
M50 241 15 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=70050 $D=1
M51 242 15 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=74680 $D=1
M52 243 241 239 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=70050 $D=1
M53 244 242 240 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=74680 $D=1
M54 237 15 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=70050 $D=1
M55 238 15 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=74680 $D=1
M56 5 16 245 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=70050 $D=1
M57 6 16 246 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=74680 $D=1
M58 247 17 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=70050 $D=1
M59 248 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=74680 $D=1
M60 249 16 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=70050 $D=1
M61 250 16 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=74680 $D=1
M62 5 249 717 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=70050 $D=1
M63 6 250 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=74680 $D=1
M64 251 717 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=70050 $D=1
M65 252 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=74680 $D=1
M66 249 245 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=70050 $D=1
M67 250 246 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=74680 $D=1
M68 251 17 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=70050 $D=1
M69 252 17 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=74680 $D=1
M70 257 18 251 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=70050 $D=1
M71 258 18 252 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=74680 $D=1
M72 255 18 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=70050 $D=1
M73 256 18 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=74680 $D=1
M74 5 19 259 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=70050 $D=1
M75 6 19 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=74680 $D=1
M76 261 20 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=70050 $D=1
M77 262 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=74680 $D=1
M78 263 19 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=70050 $D=1
M79 264 19 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=74680 $D=1
M80 5 263 719 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=70050 $D=1
M81 6 264 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=74680 $D=1
M82 265 719 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=70050 $D=1
M83 266 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=74680 $D=1
M84 263 259 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=70050 $D=1
M85 264 260 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=74680 $D=1
M86 265 20 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=70050 $D=1
M87 266 20 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=74680 $D=1
M88 257 21 265 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=70050 $D=1
M89 258 21 266 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=74680 $D=1
M90 267 21 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=70050 $D=1
M91 268 21 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=74680 $D=1
M92 5 22 269 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=70050 $D=1
M93 6 22 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=74680 $D=1
M94 271 23 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=70050 $D=1
M95 272 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=74680 $D=1
M96 273 22 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=70050 $D=1
M97 274 22 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=74680 $D=1
M98 5 273 721 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=70050 $D=1
M99 6 274 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=74680 $D=1
M100 275 721 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=70050 $D=1
M101 276 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=74680 $D=1
M102 273 269 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=70050 $D=1
M103 274 270 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=74680 $D=1
M104 275 23 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=70050 $D=1
M105 276 23 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=74680 $D=1
M106 257 24 275 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=70050 $D=1
M107 258 24 276 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=74680 $D=1
M108 277 24 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=70050 $D=1
M109 278 24 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=74680 $D=1
M110 5 25 279 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=70050 $D=1
M111 6 25 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=74680 $D=1
M112 281 26 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=70050 $D=1
M113 282 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=74680 $D=1
M114 283 25 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=70050 $D=1
M115 284 25 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=74680 $D=1
M116 5 283 723 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=70050 $D=1
M117 6 284 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=74680 $D=1
M118 285 723 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=70050 $D=1
M119 286 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=74680 $D=1
M120 283 279 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=70050 $D=1
M121 284 280 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=74680 $D=1
M122 285 26 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=70050 $D=1
M123 286 26 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=74680 $D=1
M124 257 27 285 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=70050 $D=1
M125 258 27 286 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=74680 $D=1
M126 287 27 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=70050 $D=1
M127 288 27 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=74680 $D=1
M128 5 28 289 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=70050 $D=1
M129 6 28 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=74680 $D=1
M130 291 29 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=70050 $D=1
M131 292 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=74680 $D=1
M132 293 28 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=70050 $D=1
M133 294 28 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=74680 $D=1
M134 5 293 725 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=70050 $D=1
M135 6 294 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=74680 $D=1
M136 295 725 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=70050 $D=1
M137 296 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=74680 $D=1
M138 293 289 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=70050 $D=1
M139 294 290 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=74680 $D=1
M140 295 29 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=70050 $D=1
M141 296 29 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=74680 $D=1
M142 257 30 295 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=70050 $D=1
M143 258 30 296 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=74680 $D=1
M144 297 30 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=70050 $D=1
M145 298 30 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=74680 $D=1
M146 5 31 299 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=70050 $D=1
M147 6 31 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=74680 $D=1
M148 301 32 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=70050 $D=1
M149 302 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=74680 $D=1
M150 303 31 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=70050 $D=1
M151 304 31 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=74680 $D=1
M152 5 303 727 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=70050 $D=1
M153 6 304 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=74680 $D=1
M154 305 727 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=70050 $D=1
M155 306 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=74680 $D=1
M156 303 299 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=70050 $D=1
M157 304 300 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=74680 $D=1
M158 305 32 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=70050 $D=1
M159 306 32 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=74680 $D=1
M160 257 33 305 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=70050 $D=1
M161 258 33 306 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=74680 $D=1
M162 307 33 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=70050 $D=1
M163 308 33 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=74680 $D=1
M164 5 34 309 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=70050 $D=1
M165 6 34 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=74680 $D=1
M166 311 35 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=70050 $D=1
M167 312 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=74680 $D=1
M168 313 34 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=70050 $D=1
M169 314 34 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=74680 $D=1
M170 5 313 729 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=70050 $D=1
M171 6 314 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=74680 $D=1
M172 315 729 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=70050 $D=1
M173 316 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=74680 $D=1
M174 313 309 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=70050 $D=1
M175 314 310 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=74680 $D=1
M176 315 35 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=70050 $D=1
M177 316 35 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=74680 $D=1
M178 257 36 315 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=70050 $D=1
M179 258 36 316 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=74680 $D=1
M180 317 36 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=70050 $D=1
M181 318 36 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=74680 $D=1
M182 5 37 319 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=70050 $D=1
M183 6 37 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=74680 $D=1
M184 321 38 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=70050 $D=1
M185 322 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=74680 $D=1
M186 323 37 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=70050 $D=1
M187 324 37 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=74680 $D=1
M188 5 323 731 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=70050 $D=1
M189 6 324 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=74680 $D=1
M190 325 731 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=70050 $D=1
M191 326 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=74680 $D=1
M192 323 319 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=70050 $D=1
M193 324 320 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=74680 $D=1
M194 325 38 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=70050 $D=1
M195 326 38 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=74680 $D=1
M196 257 39 325 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=70050 $D=1
M197 258 39 326 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=74680 $D=1
M198 327 39 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=70050 $D=1
M199 328 39 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=74680 $D=1
M200 5 40 329 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=70050 $D=1
M201 6 40 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=74680 $D=1
M202 331 41 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=70050 $D=1
M203 332 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=74680 $D=1
M204 333 40 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=70050 $D=1
M205 334 40 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=74680 $D=1
M206 5 333 733 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=70050 $D=1
M207 6 334 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=74680 $D=1
M208 335 733 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=70050 $D=1
M209 336 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=74680 $D=1
M210 333 329 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=70050 $D=1
M211 334 330 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=74680 $D=1
M212 335 41 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=70050 $D=1
M213 336 41 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=74680 $D=1
M214 257 42 335 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=70050 $D=1
M215 258 42 336 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=74680 $D=1
M216 337 42 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=70050 $D=1
M217 338 42 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=74680 $D=1
M218 5 43 339 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=70050 $D=1
M219 6 43 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=74680 $D=1
M220 341 44 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=70050 $D=1
M221 342 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=74680 $D=1
M222 343 43 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=70050 $D=1
M223 344 43 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=74680 $D=1
M224 5 343 735 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=70050 $D=1
M225 6 344 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=74680 $D=1
M226 345 735 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=70050 $D=1
M227 346 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=74680 $D=1
M228 343 339 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=70050 $D=1
M229 344 340 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=74680 $D=1
M230 345 44 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=70050 $D=1
M231 346 44 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=74680 $D=1
M232 257 45 345 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=70050 $D=1
M233 258 45 346 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=74680 $D=1
M234 347 45 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=70050 $D=1
M235 348 45 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=74680 $D=1
M236 5 46 349 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=70050 $D=1
M237 6 46 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=74680 $D=1
M238 351 47 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=70050 $D=1
M239 352 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=74680 $D=1
M240 353 46 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=70050 $D=1
M241 354 46 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=74680 $D=1
M242 5 353 737 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=70050 $D=1
M243 6 354 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=74680 $D=1
M244 355 737 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=70050 $D=1
M245 356 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=74680 $D=1
M246 353 349 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=70050 $D=1
M247 354 350 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=74680 $D=1
M248 355 47 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=70050 $D=1
M249 356 47 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=74680 $D=1
M250 257 48 355 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=70050 $D=1
M251 258 48 356 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=74680 $D=1
M252 357 48 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=70050 $D=1
M253 358 48 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=74680 $D=1
M254 5 49 359 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=70050 $D=1
M255 6 49 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=74680 $D=1
M256 361 50 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=70050 $D=1
M257 362 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=74680 $D=1
M258 363 49 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=70050 $D=1
M259 364 49 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=74680 $D=1
M260 5 363 739 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=70050 $D=1
M261 6 364 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=74680 $D=1
M262 365 739 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=70050 $D=1
M263 366 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=74680 $D=1
M264 363 359 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=70050 $D=1
M265 364 360 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=74680 $D=1
M266 365 50 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=70050 $D=1
M267 366 50 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=74680 $D=1
M268 257 51 365 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=70050 $D=1
M269 258 51 366 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=74680 $D=1
M270 367 51 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=70050 $D=1
M271 368 51 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=74680 $D=1
M272 5 52 369 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=70050 $D=1
M273 6 52 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=74680 $D=1
M274 371 53 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=70050 $D=1
M275 372 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=74680 $D=1
M276 373 52 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=70050 $D=1
M277 374 52 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=74680 $D=1
M278 5 373 741 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=70050 $D=1
M279 6 374 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=74680 $D=1
M280 375 741 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=70050 $D=1
M281 376 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=74680 $D=1
M282 373 369 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=70050 $D=1
M283 374 370 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=74680 $D=1
M284 375 53 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=70050 $D=1
M285 376 53 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=74680 $D=1
M286 257 54 375 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=70050 $D=1
M287 258 54 376 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=74680 $D=1
M288 377 54 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=70050 $D=1
M289 378 54 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=74680 $D=1
M290 5 55 379 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=70050 $D=1
M291 6 55 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=74680 $D=1
M292 381 56 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=70050 $D=1
M293 382 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=74680 $D=1
M294 383 55 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=70050 $D=1
M295 384 55 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=74680 $D=1
M296 5 383 743 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=70050 $D=1
M297 6 384 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=74680 $D=1
M298 385 743 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=70050 $D=1
M299 386 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=74680 $D=1
M300 383 379 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=70050 $D=1
M301 384 380 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=74680 $D=1
M302 385 56 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=70050 $D=1
M303 386 56 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=74680 $D=1
M304 257 57 385 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=70050 $D=1
M305 258 57 386 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=74680 $D=1
M306 387 57 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=70050 $D=1
M307 388 57 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=74680 $D=1
M308 5 58 389 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=70050 $D=1
M309 6 58 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=74680 $D=1
M310 391 59 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=70050 $D=1
M311 392 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=74680 $D=1
M312 393 58 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=70050 $D=1
M313 394 58 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=74680 $D=1
M314 5 393 745 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=70050 $D=1
M315 6 394 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=74680 $D=1
M316 395 745 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=70050 $D=1
M317 396 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=74680 $D=1
M318 393 389 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=70050 $D=1
M319 394 390 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=74680 $D=1
M320 395 59 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=70050 $D=1
M321 396 59 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=74680 $D=1
M322 257 60 395 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=70050 $D=1
M323 258 60 396 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=74680 $D=1
M324 397 60 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=70050 $D=1
M325 398 60 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=74680 $D=1
M326 5 61 399 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=70050 $D=1
M327 6 61 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=74680 $D=1
M328 401 62 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=70050 $D=1
M329 402 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=74680 $D=1
M330 403 61 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=70050 $D=1
M331 404 61 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=74680 $D=1
M332 5 403 747 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=70050 $D=1
M333 6 404 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=74680 $D=1
M334 405 747 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=70050 $D=1
M335 406 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=74680 $D=1
M336 403 399 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=70050 $D=1
M337 404 400 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=74680 $D=1
M338 405 62 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=70050 $D=1
M339 406 62 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=74680 $D=1
M340 257 63 405 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=70050 $D=1
M341 258 63 406 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=74680 $D=1
M342 407 63 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=70050 $D=1
M343 408 63 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=74680 $D=1
M344 5 64 409 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=70050 $D=1
M345 6 64 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=74680 $D=1
M346 411 65 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=70050 $D=1
M347 412 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=74680 $D=1
M348 413 64 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=70050 $D=1
M349 414 64 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=74680 $D=1
M350 5 413 749 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=70050 $D=1
M351 6 414 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=74680 $D=1
M352 415 749 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=70050 $D=1
M353 416 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=74680 $D=1
M354 413 409 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=70050 $D=1
M355 414 410 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=74680 $D=1
M356 415 65 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=70050 $D=1
M357 416 65 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=74680 $D=1
M358 257 66 415 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=70050 $D=1
M359 258 66 416 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=74680 $D=1
M360 417 66 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=70050 $D=1
M361 418 66 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=74680 $D=1
M362 5 67 419 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=70050 $D=1
M363 6 67 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=74680 $D=1
M364 421 68 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=70050 $D=1
M365 422 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=74680 $D=1
M366 423 67 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=70050 $D=1
M367 424 67 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=74680 $D=1
M368 5 423 751 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=70050 $D=1
M369 6 424 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=74680 $D=1
M370 425 751 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=70050 $D=1
M371 426 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=74680 $D=1
M372 423 419 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=70050 $D=1
M373 424 420 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=74680 $D=1
M374 425 68 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=70050 $D=1
M375 426 68 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=74680 $D=1
M376 257 69 425 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=70050 $D=1
M377 258 69 426 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=74680 $D=1
M378 427 69 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=70050 $D=1
M379 428 69 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=74680 $D=1
M380 5 70 429 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=70050 $D=1
M381 6 70 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=74680 $D=1
M382 431 71 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=70050 $D=1
M383 432 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=74680 $D=1
M384 433 70 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=70050 $D=1
M385 434 70 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=74680 $D=1
M386 5 433 753 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=70050 $D=1
M387 6 434 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=74680 $D=1
M388 435 753 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=70050 $D=1
M389 436 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=74680 $D=1
M390 433 429 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=70050 $D=1
M391 434 430 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=74680 $D=1
M392 435 71 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=70050 $D=1
M393 436 71 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=74680 $D=1
M394 257 72 435 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=70050 $D=1
M395 258 72 436 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=74680 $D=1
M396 437 72 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=70050 $D=1
M397 438 72 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=74680 $D=1
M398 5 73 439 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=70050 $D=1
M399 6 73 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=74680 $D=1
M400 441 74 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=70050 $D=1
M401 442 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=74680 $D=1
M402 443 73 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=70050 $D=1
M403 444 73 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=74680 $D=1
M404 5 443 755 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=70050 $D=1
M405 6 444 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=74680 $D=1
M406 445 755 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=70050 $D=1
M407 446 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=74680 $D=1
M408 443 439 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=70050 $D=1
M409 444 440 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=74680 $D=1
M410 445 74 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=70050 $D=1
M411 446 74 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=74680 $D=1
M412 257 75 445 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=70050 $D=1
M413 258 75 446 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=74680 $D=1
M414 447 75 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=70050 $D=1
M415 448 75 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=74680 $D=1
M416 5 76 449 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=70050 $D=1
M417 6 76 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=74680 $D=1
M418 451 77 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=70050 $D=1
M419 452 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=74680 $D=1
M420 453 76 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=70050 $D=1
M421 454 76 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=74680 $D=1
M422 5 453 757 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=70050 $D=1
M423 6 454 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=74680 $D=1
M424 455 757 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=70050 $D=1
M425 456 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=74680 $D=1
M426 453 449 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=70050 $D=1
M427 454 450 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=74680 $D=1
M428 455 77 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=70050 $D=1
M429 456 77 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=74680 $D=1
M430 257 78 455 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=70050 $D=1
M431 258 78 456 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=74680 $D=1
M432 457 78 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=70050 $D=1
M433 458 78 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=74680 $D=1
M434 5 79 459 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=70050 $D=1
M435 6 79 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=74680 $D=1
M436 461 80 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=70050 $D=1
M437 462 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=74680 $D=1
M438 463 79 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=70050 $D=1
M439 464 79 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=74680 $D=1
M440 5 463 759 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=70050 $D=1
M441 6 464 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=74680 $D=1
M442 465 759 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=70050 $D=1
M443 466 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=74680 $D=1
M444 463 459 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=70050 $D=1
M445 464 460 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=74680 $D=1
M446 465 80 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=70050 $D=1
M447 466 80 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=74680 $D=1
M448 257 81 465 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=70050 $D=1
M449 258 81 466 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=74680 $D=1
M450 467 81 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=70050 $D=1
M451 468 81 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=74680 $D=1
M452 5 82 469 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=70050 $D=1
M453 6 82 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=74680 $D=1
M454 471 83 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=70050 $D=1
M455 472 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=74680 $D=1
M456 473 82 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=70050 $D=1
M457 474 82 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=74680 $D=1
M458 5 473 761 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=70050 $D=1
M459 6 474 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=74680 $D=1
M460 475 761 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=70050 $D=1
M461 476 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=74680 $D=1
M462 473 469 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=70050 $D=1
M463 474 470 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=74680 $D=1
M464 475 83 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=70050 $D=1
M465 476 83 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=74680 $D=1
M466 257 84 475 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=70050 $D=1
M467 258 84 476 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=74680 $D=1
M468 477 84 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=70050 $D=1
M469 478 84 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=74680 $D=1
M470 5 85 479 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=70050 $D=1
M471 6 85 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=74680 $D=1
M472 481 86 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=70050 $D=1
M473 482 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=74680 $D=1
M474 483 85 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=70050 $D=1
M475 484 85 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=74680 $D=1
M476 5 483 763 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=70050 $D=1
M477 6 484 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=74680 $D=1
M478 485 763 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=70050 $D=1
M479 486 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=74680 $D=1
M480 483 479 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=70050 $D=1
M481 484 480 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=74680 $D=1
M482 485 86 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=70050 $D=1
M483 486 86 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=74680 $D=1
M484 257 87 485 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=70050 $D=1
M485 258 87 486 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=74680 $D=1
M486 487 87 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=70050 $D=1
M487 488 87 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=74680 $D=1
M488 5 88 489 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=70050 $D=1
M489 6 88 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=74680 $D=1
M490 491 89 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=70050 $D=1
M491 492 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=74680 $D=1
M492 493 88 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=70050 $D=1
M493 494 88 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=74680 $D=1
M494 5 493 765 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=70050 $D=1
M495 6 494 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=74680 $D=1
M496 495 765 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=70050 $D=1
M497 496 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=74680 $D=1
M498 493 489 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=70050 $D=1
M499 494 490 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=74680 $D=1
M500 495 89 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=70050 $D=1
M501 496 89 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=74680 $D=1
M502 257 90 495 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=70050 $D=1
M503 258 90 496 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=74680 $D=1
M504 497 90 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=70050 $D=1
M505 498 90 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=74680 $D=1
M506 5 91 499 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=70050 $D=1
M507 6 91 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=74680 $D=1
M508 501 92 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=70050 $D=1
M509 502 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=74680 $D=1
M510 503 91 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=70050 $D=1
M511 504 91 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=74680 $D=1
M512 5 503 767 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=70050 $D=1
M513 6 504 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=74680 $D=1
M514 505 767 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=70050 $D=1
M515 506 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=74680 $D=1
M516 503 499 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=70050 $D=1
M517 504 500 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=74680 $D=1
M518 505 92 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=70050 $D=1
M519 506 92 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=74680 $D=1
M520 257 93 505 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=70050 $D=1
M521 258 93 506 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=74680 $D=1
M522 507 93 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=70050 $D=1
M523 508 93 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=74680 $D=1
M524 5 94 509 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=70050 $D=1
M525 6 94 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=74680 $D=1
M526 511 95 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=70050 $D=1
M527 512 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=74680 $D=1
M528 513 94 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=70050 $D=1
M529 514 94 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=74680 $D=1
M530 5 513 769 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=70050 $D=1
M531 6 514 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=74680 $D=1
M532 515 769 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=70050 $D=1
M533 516 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=74680 $D=1
M534 513 509 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=70050 $D=1
M535 514 510 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=74680 $D=1
M536 515 95 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=70050 $D=1
M537 516 95 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=74680 $D=1
M538 257 96 515 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=70050 $D=1
M539 258 96 516 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=74680 $D=1
M540 517 96 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=70050 $D=1
M541 518 96 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=74680 $D=1
M542 5 97 519 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=70050 $D=1
M543 6 97 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=74680 $D=1
M544 521 98 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=70050 $D=1
M545 522 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=74680 $D=1
M546 523 97 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=70050 $D=1
M547 524 97 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=74680 $D=1
M548 5 523 771 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=70050 $D=1
M549 6 524 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=74680 $D=1
M550 525 771 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=70050 $D=1
M551 526 772 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=74680 $D=1
M552 523 519 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=70050 $D=1
M553 524 520 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=74680 $D=1
M554 525 98 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=70050 $D=1
M555 526 98 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=74680 $D=1
M556 257 99 525 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=70050 $D=1
M557 258 99 526 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=74680 $D=1
M558 527 99 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=70050 $D=1
M559 528 99 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=74680 $D=1
M560 5 100 529 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=70050 $D=1
M561 6 100 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=74680 $D=1
M562 531 101 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=70050 $D=1
M563 532 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=74680 $D=1
M564 533 100 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=70050 $D=1
M565 534 100 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=74680 $D=1
M566 5 533 773 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=70050 $D=1
M567 6 534 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=74680 $D=1
M568 535 773 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=70050 $D=1
M569 536 774 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=74680 $D=1
M570 533 529 535 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=70050 $D=1
M571 534 530 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=74680 $D=1
M572 535 101 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=70050 $D=1
M573 536 101 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=74680 $D=1
M574 257 102 535 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=70050 $D=1
M575 258 102 536 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=74680 $D=1
M576 537 102 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=70050 $D=1
M577 538 102 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=74680 $D=1
M578 5 103 539 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=70050 $D=1
M579 6 103 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=74680 $D=1
M580 541 104 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=70050 $D=1
M581 542 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=74680 $D=1
M582 543 103 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=70050 $D=1
M583 544 103 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=74680 $D=1
M584 5 543 775 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=70050 $D=1
M585 6 544 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=74680 $D=1
M586 545 775 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=70050 $D=1
M587 546 776 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=74680 $D=1
M588 543 539 545 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=70050 $D=1
M589 544 540 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=74680 $D=1
M590 545 104 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=70050 $D=1
M591 546 104 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=74680 $D=1
M592 257 105 545 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=70050 $D=1
M593 258 105 546 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=74680 $D=1
M594 547 105 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=70050 $D=1
M595 548 105 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=74680 $D=1
M596 5 106 549 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=70050 $D=1
M597 6 106 550 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=74680 $D=1
M598 551 107 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=70050 $D=1
M599 552 107 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=74680 $D=1
M600 553 106 243 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=70050 $D=1
M601 554 106 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=74680 $D=1
M602 5 553 777 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=70050 $D=1
M603 6 554 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=74680 $D=1
M604 555 777 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=70050 $D=1
M605 556 778 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=74680 $D=1
M606 553 549 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=70050 $D=1
M607 554 550 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=74680 $D=1
M608 555 107 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=70050 $D=1
M609 556 107 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=74680 $D=1
M610 257 109 555 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=70050 $D=1
M611 258 109 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=74680 $D=1
M612 557 109 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=70050 $D=1
M613 558 109 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=74680 $D=1
M614 5 110 559 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=70050 $D=1
M615 6 110 560 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=74680 $D=1
M616 561 111 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=70050 $D=1
M617 562 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=74680 $D=1
M618 5 111 253 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=70050 $D=1
M619 6 111 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=74680 $D=1
M620 257 110 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=70050 $D=1
M621 258 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=74680 $D=1
M622 5 565 563 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=70050 $D=1
M623 6 566 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=74680 $D=1
M624 565 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=70050 $D=1
M625 566 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=74680 $D=1
M626 779 253 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=70050 $D=1
M627 780 254 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=74680 $D=1
M628 567 563 779 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=70050 $D=1
M629 568 564 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=74680 $D=1
M630 5 567 569 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=70050 $D=1
M631 6 568 570 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=74680 $D=1
M632 781 569 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=70050 $D=1
M633 782 570 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=74680 $D=1
M634 567 565 781 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=70050 $D=1
M635 568 566 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=74680 $D=1
M636 5 573 571 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=70050 $D=1
M637 6 574 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=74680 $D=1
M638 573 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=70050 $D=1
M639 574 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=74680 $D=1
M640 783 257 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=70050 $D=1
M641 784 258 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=74680 $D=1
M642 575 571 783 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=70050 $D=1
M643 576 572 784 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=74680 $D=1
M644 5 575 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=70050 $D=1
M645 6 576 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=74680 $D=1
M646 785 116 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=70050 $D=1
M647 786 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=74680 $D=1
M648 575 573 785 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=70050 $D=1
M649 576 574 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=74680 $D=1
M650 577 120 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=70050 $D=1
M651 578 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=74680 $D=1
M652 579 577 569 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=70050 $D=1
M653 580 578 570 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=74680 $D=1
M654 121 120 579 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=70050 $D=1
M655 121 120 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=74680 $D=1
M656 581 122 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=70050 $D=1
M657 582 122 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=74680 $D=1
M658 583 581 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=70050 $D=1
M659 584 582 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=74680 $D=1
M660 787 122 583 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=70050 $D=1
M661 788 122 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=74680 $D=1
M662 5 116 787 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=70050 $D=1
M663 6 117 788 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=74680 $D=1
M664 585 123 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=70050 $D=1
M665 586 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=74680 $D=1
M666 587 585 583 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=70050 $D=1
M667 588 586 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=74680 $D=1
M668 10 123 587 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=70050 $D=1
M669 11 123 588 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=74680 $D=1
M670 590 589 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=70050 $D=1
M671 591 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=74680 $D=1
M672 5 594 592 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=70050 $D=1
M673 6 595 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=74680 $D=1
M674 596 579 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=70050 $D=1
M675 597 580 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=74680 $D=1
M676 594 596 589 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=70050 $D=1
M677 595 597 124 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=74680 $D=1
M678 590 579 594 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=70050 $D=1
M679 591 580 595 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=74680 $D=1
M680 598 592 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=70050 $D=1
M681 599 593 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=74680 $D=1
M682 125 598 587 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=70050 $D=1
M683 589 599 588 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=74680 $D=1
M684 579 592 125 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=70050 $D=1
M685 580 593 589 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=74680 $D=1
M686 600 125 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=70050 $D=1
M687 601 589 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=74680 $D=1
M688 602 592 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=70050 $D=1
M689 603 593 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=74680 $D=1
M690 604 602 600 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=70050 $D=1
M691 605 603 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=74680 $D=1
M692 587 592 604 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=70050 $D=1
M693 588 593 605 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=74680 $D=1
M694 606 579 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=70050 $D=1
M695 607 580 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=74680 $D=1
M696 5 587 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=70050 $D=1
M697 6 588 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=74680 $D=1
M698 608 604 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=70050 $D=1
M699 609 605 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=74680 $D=1
M700 807 579 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=70050 $D=1
M701 808 580 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=74680 $D=1
M702 610 587 807 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=70050 $D=1
M703 611 588 808 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=74680 $D=1
M704 809 579 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=70050 $D=1
M705 810 580 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=74680 $D=1
M706 612 587 809 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=70050 $D=1
M707 613 588 810 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=74680 $D=1
M708 616 579 614 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=70050 $D=1
M709 617 580 615 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=74680 $D=1
M710 614 587 616 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=70050 $D=1
M711 615 588 617 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=74680 $D=1
M712 5 612 614 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=70050 $D=1
M713 6 613 615 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=74680 $D=1
M714 618 128 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=70050 $D=1
M715 619 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=74680 $D=1
M716 620 618 606 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=70050 $D=1
M717 621 619 607 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=74680 $D=1
M718 610 128 620 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=70050 $D=1
M719 611 128 621 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=74680 $D=1
M720 622 618 608 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=70050 $D=1
M721 623 619 609 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=74680 $D=1
M722 616 128 622 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=70050 $D=1
M723 617 128 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=74680 $D=1
M724 624 129 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=70050 $D=1
M725 625 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=74680 $D=1
M726 626 624 622 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=70050 $D=1
M727 627 625 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=74680 $D=1
M728 620 129 626 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=70050 $D=1
M729 621 129 627 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=74680 $D=1
M730 12 626 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=70050 $D=1
M731 13 627 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=74680 $D=1
M732 628 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=70050 $D=1
M733 629 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=74680 $D=1
M734 630 628 131 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=70050 $D=1
M735 631 629 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=74680 $D=1
M736 133 130 630 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=70050 $D=1
M737 134 130 631 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=74680 $D=1
M738 632 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=70050 $D=1
M739 633 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=74680 $D=1
M740 634 632 135 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=70050 $D=1
M741 635 633 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=74680 $D=1
M742 137 130 634 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=70050 $D=1
M743 138 130 635 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=74680 $D=1
M744 636 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=70050 $D=1
M745 637 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=74680 $D=1
M746 638 636 126 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=70050 $D=1
M747 639 637 139 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=74680 $D=1
M748 114 130 638 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=70050 $D=1
M749 115 130 639 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=74680 $D=1
M750 640 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=70050 $D=1
M751 641 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=74680 $D=1
M752 642 640 140 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=70050 $D=1
M753 643 641 141 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=74680 $D=1
M754 142 130 642 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=70050 $D=1
M755 143 130 643 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=74680 $D=1
M756 644 130 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=70050 $D=1
M757 645 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=74680 $D=1
M758 646 644 144 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=70050 $D=1
M759 647 645 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=74680 $D=1
M760 145 130 646 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=70050 $D=1
M761 146 130 647 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=74680 $D=1
M762 5 579 789 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=70050 $D=1
M763 6 580 790 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=74680 $D=1
M764 134 789 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=70050 $D=1
M765 131 790 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=74680 $D=1
M766 648 147 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=70050 $D=1
M767 649 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=74680 $D=1
M768 149 648 134 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=70050 $D=1
M769 150 649 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=74680 $D=1
M770 630 147 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=70050 $D=1
M771 631 147 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=74680 $D=1
M772 650 151 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=70050 $D=1
M773 651 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=74680 $D=1
M774 118 650 149 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=70050 $D=1
M775 119 651 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=74680 $D=1
M776 634 151 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=70050 $D=1
M777 635 151 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=74680 $D=1
M778 652 152 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=70050 $D=1
M779 653 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=74680 $D=1
M780 108 652 118 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=70050 $D=1
M781 113 653 119 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=74680 $D=1
M782 638 152 108 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=70050 $D=1
M783 639 152 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=74680 $D=1
M784 654 153 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=70050 $D=1
M785 655 153 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=74680 $D=1
M786 148 654 108 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=70050 $D=1
M787 154 655 113 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=74680 $D=1
M788 642 153 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=70050 $D=1
M789 643 153 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=74680 $D=1
M790 656 155 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=70050 $D=1
M791 657 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=74680 $D=1
M792 229 656 148 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=70050 $D=1
M793 230 657 154 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=74680 $D=1
M794 646 155 229 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=70050 $D=1
M795 647 155 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=74680 $D=1
M796 658 156 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=70050 $D=1
M797 659 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=74680 $D=1
M798 660 658 116 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=70050 $D=1
M799 661 659 117 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=74680 $D=1
M800 10 156 660 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=70050 $D=1
M801 11 156 661 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=74680 $D=1
M802 811 569 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=70050 $D=1
M803 812 570 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=74680 $D=1
M804 662 660 811 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=70050 $D=1
M805 663 661 812 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=74680 $D=1
M806 666 569 664 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=70050 $D=1
M807 667 570 665 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=74680 $D=1
M808 664 660 666 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=70050 $D=1
M809 665 661 667 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=74680 $D=1
M810 5 662 664 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=70050 $D=1
M811 6 663 665 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=74680 $D=1
M812 813 157 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=70050 $D=1
M813 814 668 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=74680 $D=1
M814 791 666 813 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=70050 $D=1
M815 792 667 814 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=74680 $D=1
M816 668 791 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=70050 $D=1
M817 158 792 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=74680 $D=1
M818 669 569 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=70050 $D=1
M819 670 570 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=74680 $D=1
M820 5 671 669 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=70050 $D=1
M821 6 672 670 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=74680 $D=1
M822 671 660 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=70050 $D=1
M823 672 661 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=74680 $D=1
M824 815 669 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=70050 $D=1
M825 816 670 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=74680 $D=1
M826 673 157 815 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=70050 $D=1
M827 674 668 816 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=74680 $D=1
M828 676 159 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=70050 $D=1
M829 677 675 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=74680 $D=1
M830 817 673 5 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=70050 $D=1
M831 818 674 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=74680 $D=1
M832 675 676 817 5 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=70050 $D=1
M833 160 677 818 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=74680 $D=1
M834 679 678 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=70050 $D=1
M835 680 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=74680 $D=1
M836 5 683 681 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=70050 $D=1
M837 6 684 682 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=74680 $D=1
M838 685 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=70050 $D=1
M839 686 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=74680 $D=1
M840 683 685 678 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=70050 $D=1
M841 684 686 161 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=74680 $D=1
M842 679 121 683 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=70050 $D=1
M843 680 121 684 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=74680 $D=1
M844 687 681 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=70050 $D=1
M845 688 682 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=74680 $D=1
M846 162 687 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=70050 $D=1
M847 678 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=74680 $D=1
M848 121 681 162 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=70050 $D=1
M849 121 682 678 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=74680 $D=1
M850 689 162 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=70050 $D=1
M851 690 678 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=74680 $D=1
M852 691 681 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=70050 $D=1
M853 692 682 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=74680 $D=1
M854 231 691 689 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=70050 $D=1
M855 232 692 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=74680 $D=1
M856 5 681 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=70050 $D=1
M857 6 682 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=74680 $D=1
M858 693 163 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=70050 $D=1
M859 694 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=74680 $D=1
M860 695 693 231 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=70050 $D=1
M861 696 694 232 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=74680 $D=1
M862 12 163 695 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=70050 $D=1
M863 13 163 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=74680 $D=1
M864 697 164 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=70050 $D=1
M865 698 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=74680 $D=1
M866 164 697 695 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=70050 $D=1
M867 164 698 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=74680 $D=1
M868 5 164 164 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=70050 $D=1
M869 6 164 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=74680 $D=1
M870 699 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=70050 $D=1
M871 700 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=74680 $D=1
M872 5 699 701 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=70050 $D=1
M873 6 700 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=74680 $D=1
M874 703 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=70050 $D=1
M875 704 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=74680 $D=1
M876 705 699 164 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=70050 $D=1
M877 706 700 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=74680 $D=1
M878 5 705 793 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=70050 $D=1
M879 6 706 794 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=74680 $D=1
M880 707 793 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=70050 $D=1
M881 708 794 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=74680 $D=1
M882 705 701 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=70050 $D=1
M883 706 702 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=74680 $D=1
M884 709 112 707 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=70050 $D=1
M885 710 112 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=74680 $D=1
M886 5 713 711 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=70050 $D=1
M887 6 714 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=74680 $D=1
M888 713 112 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=70050 $D=1
M889 714 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=74680 $D=1
M890 795 709 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=70050 $D=1
M891 796 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=74680 $D=1
M892 715 711 795 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=70050 $D=1
M893 716 712 796 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=74680 $D=1
M894 5 715 121 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=70050 $D=1
M895 6 716 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=74680 $D=1
M896 797 121 5 5 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=70050 $D=1
M897 798 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=74680 $D=1
M898 715 713 797 5 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=70050 $D=1
M899 716 714 798 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=74680 $D=1
M900 205 1 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=71300 $D=0
M901 206 1 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=75930 $D=0
M902 207 1 2 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=71300 $D=0
M903 208 1 3 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=75930 $D=0
M904 5 205 207 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=71300 $D=0
M905 6 206 208 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=75930 $D=0
M906 209 1 4 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=71300 $D=0
M907 210 1 4 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=75930 $D=0
M908 3 205 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=71300 $D=0
M909 3 206 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=75930 $D=0
M910 211 1 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=71300 $D=0
M911 212 1 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=75930 $D=0
M912 5 205 211 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=71300 $D=0
M913 3 206 212 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=75930 $D=0
M914 215 7 211 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=71300 $D=0
M915 216 7 212 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=75930 $D=0
M916 213 7 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=71300 $D=0
M917 214 7 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=75930 $D=0
M918 217 7 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=71300 $D=0
M919 218 7 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=75930 $D=0
M920 207 213 217 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=71300 $D=0
M921 208 214 218 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=75930 $D=0
M922 219 8 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=71300 $D=0
M923 220 8 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=75930 $D=0
M924 221 8 217 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=71300 $D=0
M925 222 8 218 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=75930 $D=0
M926 215 219 221 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=71300 $D=0
M927 216 220 222 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=75930 $D=0
M928 223 9 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=71300 $D=0
M929 224 9 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=75930 $D=0
M930 225 9 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=71300 $D=0
M931 226 9 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=75930 $D=0
M932 10 223 225 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=71300 $D=0
M933 11 224 226 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=75930 $D=0
M934 227 9 12 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=71300 $D=0
M935 228 9 13 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=75930 $D=0
M936 229 223 227 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=71300 $D=0
M937 230 224 228 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=75930 $D=0
M938 233 9 231 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=71300 $D=0
M939 234 9 232 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=75930 $D=0
M940 221 223 233 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=71300 $D=0
M941 222 224 234 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=75930 $D=0
M942 237 14 233 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=71300 $D=0
M943 238 14 234 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=75930 $D=0
M944 235 14 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=71300 $D=0
M945 236 14 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=75930 $D=0
M946 239 14 227 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=71300 $D=0
M947 240 14 228 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=75930 $D=0
M948 225 235 239 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=71300 $D=0
M949 226 236 240 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=75930 $D=0
M950 241 15 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=71300 $D=0
M951 242 15 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=75930 $D=0
M952 243 15 239 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=71300 $D=0
M953 244 15 240 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=75930 $D=0
M954 237 241 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=71300 $D=0
M955 238 242 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=75930 $D=0
M956 165 16 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=71300 $D=0
M957 166 16 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=75930 $D=0
M958 247 17 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=71300 $D=0
M959 248 17 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=75930 $D=0
M960 249 245 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=71300 $D=0
M961 250 246 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=75930 $D=0
M962 165 249 717 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=71300 $D=0
M963 166 250 718 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=75930 $D=0
M964 251 717 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=71300 $D=0
M965 252 718 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=75930 $D=0
M966 249 16 251 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=71300 $D=0
M967 250 16 252 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=75930 $D=0
M968 251 247 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=71300 $D=0
M969 252 248 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=75930 $D=0
M970 257 255 251 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=71300 $D=0
M971 258 256 252 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=75930 $D=0
M972 255 18 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=71300 $D=0
M973 256 18 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=75930 $D=0
M974 165 19 259 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=71300 $D=0
M975 166 19 260 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=75930 $D=0
M976 261 20 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=71300 $D=0
M977 262 20 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=75930 $D=0
M978 263 259 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=71300 $D=0
M979 264 260 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=75930 $D=0
M980 165 263 719 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=71300 $D=0
M981 166 264 720 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=75930 $D=0
M982 265 719 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=71300 $D=0
M983 266 720 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=75930 $D=0
M984 263 19 265 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=71300 $D=0
M985 264 19 266 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=75930 $D=0
M986 265 261 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=71300 $D=0
M987 266 262 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=75930 $D=0
M988 257 267 265 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=71300 $D=0
M989 258 268 266 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=75930 $D=0
M990 267 21 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=71300 $D=0
M991 268 21 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=75930 $D=0
M992 165 22 269 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=71300 $D=0
M993 166 22 270 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=75930 $D=0
M994 271 23 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=71300 $D=0
M995 272 23 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=75930 $D=0
M996 273 269 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=71300 $D=0
M997 274 270 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=75930 $D=0
M998 165 273 721 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=71300 $D=0
M999 166 274 722 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=75930 $D=0
M1000 275 721 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=71300 $D=0
M1001 276 722 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=75930 $D=0
M1002 273 22 275 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=71300 $D=0
M1003 274 22 276 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=75930 $D=0
M1004 275 271 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=71300 $D=0
M1005 276 272 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=75930 $D=0
M1006 257 277 275 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=71300 $D=0
M1007 258 278 276 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=75930 $D=0
M1008 277 24 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=71300 $D=0
M1009 278 24 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=75930 $D=0
M1010 165 25 279 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=71300 $D=0
M1011 166 25 280 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=75930 $D=0
M1012 281 26 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=71300 $D=0
M1013 282 26 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=75930 $D=0
M1014 283 279 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=71300 $D=0
M1015 284 280 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=75930 $D=0
M1016 165 283 723 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=71300 $D=0
M1017 166 284 724 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=75930 $D=0
M1018 285 723 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=71300 $D=0
M1019 286 724 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=75930 $D=0
M1020 283 25 285 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=71300 $D=0
M1021 284 25 286 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=75930 $D=0
M1022 285 281 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=71300 $D=0
M1023 286 282 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=75930 $D=0
M1024 257 287 285 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=71300 $D=0
M1025 258 288 286 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=75930 $D=0
M1026 287 27 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=71300 $D=0
M1027 288 27 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=75930 $D=0
M1028 165 28 289 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=71300 $D=0
M1029 166 28 290 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=75930 $D=0
M1030 291 29 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=71300 $D=0
M1031 292 29 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=75930 $D=0
M1032 293 289 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=71300 $D=0
M1033 294 290 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=75930 $D=0
M1034 165 293 725 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=71300 $D=0
M1035 166 294 726 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=75930 $D=0
M1036 295 725 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=71300 $D=0
M1037 296 726 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=75930 $D=0
M1038 293 28 295 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=71300 $D=0
M1039 294 28 296 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=75930 $D=0
M1040 295 291 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=71300 $D=0
M1041 296 292 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=75930 $D=0
M1042 257 297 295 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=71300 $D=0
M1043 258 298 296 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=75930 $D=0
M1044 297 30 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=71300 $D=0
M1045 298 30 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=75930 $D=0
M1046 165 31 299 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=71300 $D=0
M1047 166 31 300 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=75930 $D=0
M1048 301 32 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=71300 $D=0
M1049 302 32 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=75930 $D=0
M1050 303 299 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=71300 $D=0
M1051 304 300 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=75930 $D=0
M1052 165 303 727 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=71300 $D=0
M1053 166 304 728 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=75930 $D=0
M1054 305 727 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=71300 $D=0
M1055 306 728 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=75930 $D=0
M1056 303 31 305 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=71300 $D=0
M1057 304 31 306 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=75930 $D=0
M1058 305 301 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=71300 $D=0
M1059 306 302 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=75930 $D=0
M1060 257 307 305 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=71300 $D=0
M1061 258 308 306 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=75930 $D=0
M1062 307 33 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=71300 $D=0
M1063 308 33 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=75930 $D=0
M1064 165 34 309 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=71300 $D=0
M1065 166 34 310 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=75930 $D=0
M1066 311 35 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=71300 $D=0
M1067 312 35 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=75930 $D=0
M1068 313 309 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=71300 $D=0
M1069 314 310 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=75930 $D=0
M1070 165 313 729 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=71300 $D=0
M1071 166 314 730 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=75930 $D=0
M1072 315 729 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=71300 $D=0
M1073 316 730 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=75930 $D=0
M1074 313 34 315 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=71300 $D=0
M1075 314 34 316 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=75930 $D=0
M1076 315 311 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=71300 $D=0
M1077 316 312 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=75930 $D=0
M1078 257 317 315 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=71300 $D=0
M1079 258 318 316 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=75930 $D=0
M1080 317 36 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=71300 $D=0
M1081 318 36 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=75930 $D=0
M1082 165 37 319 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=71300 $D=0
M1083 166 37 320 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=75930 $D=0
M1084 321 38 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=71300 $D=0
M1085 322 38 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=75930 $D=0
M1086 323 319 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=71300 $D=0
M1087 324 320 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=75930 $D=0
M1088 165 323 731 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=71300 $D=0
M1089 166 324 732 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=75930 $D=0
M1090 325 731 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=71300 $D=0
M1091 326 732 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=75930 $D=0
M1092 323 37 325 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=71300 $D=0
M1093 324 37 326 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=75930 $D=0
M1094 325 321 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=71300 $D=0
M1095 326 322 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=75930 $D=0
M1096 257 327 325 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=71300 $D=0
M1097 258 328 326 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=75930 $D=0
M1098 327 39 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=71300 $D=0
M1099 328 39 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=75930 $D=0
M1100 165 40 329 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=71300 $D=0
M1101 166 40 330 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=75930 $D=0
M1102 331 41 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=71300 $D=0
M1103 332 41 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=75930 $D=0
M1104 333 329 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=71300 $D=0
M1105 334 330 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=75930 $D=0
M1106 165 333 733 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=71300 $D=0
M1107 166 334 734 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=75930 $D=0
M1108 335 733 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=71300 $D=0
M1109 336 734 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=75930 $D=0
M1110 333 40 335 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=71300 $D=0
M1111 334 40 336 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=75930 $D=0
M1112 335 331 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=71300 $D=0
M1113 336 332 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=75930 $D=0
M1114 257 337 335 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=71300 $D=0
M1115 258 338 336 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=75930 $D=0
M1116 337 42 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=71300 $D=0
M1117 338 42 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=75930 $D=0
M1118 165 43 339 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=71300 $D=0
M1119 166 43 340 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=75930 $D=0
M1120 341 44 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=71300 $D=0
M1121 342 44 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=75930 $D=0
M1122 343 339 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=71300 $D=0
M1123 344 340 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=75930 $D=0
M1124 165 343 735 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=71300 $D=0
M1125 166 344 736 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=75930 $D=0
M1126 345 735 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=71300 $D=0
M1127 346 736 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=75930 $D=0
M1128 343 43 345 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=71300 $D=0
M1129 344 43 346 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=75930 $D=0
M1130 345 341 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=71300 $D=0
M1131 346 342 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=75930 $D=0
M1132 257 347 345 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=71300 $D=0
M1133 258 348 346 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=75930 $D=0
M1134 347 45 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=71300 $D=0
M1135 348 45 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=75930 $D=0
M1136 165 46 349 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=71300 $D=0
M1137 166 46 350 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=75930 $D=0
M1138 351 47 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=71300 $D=0
M1139 352 47 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=75930 $D=0
M1140 353 349 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=71300 $D=0
M1141 354 350 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=75930 $D=0
M1142 165 353 737 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=71300 $D=0
M1143 166 354 738 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=75930 $D=0
M1144 355 737 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=71300 $D=0
M1145 356 738 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=75930 $D=0
M1146 353 46 355 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=71300 $D=0
M1147 354 46 356 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=75930 $D=0
M1148 355 351 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=71300 $D=0
M1149 356 352 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=75930 $D=0
M1150 257 357 355 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=71300 $D=0
M1151 258 358 356 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=75930 $D=0
M1152 357 48 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=71300 $D=0
M1153 358 48 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=75930 $D=0
M1154 165 49 359 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=71300 $D=0
M1155 166 49 360 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=75930 $D=0
M1156 361 50 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=71300 $D=0
M1157 362 50 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=75930 $D=0
M1158 363 359 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=71300 $D=0
M1159 364 360 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=75930 $D=0
M1160 165 363 739 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=71300 $D=0
M1161 166 364 740 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=75930 $D=0
M1162 365 739 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=71300 $D=0
M1163 366 740 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=75930 $D=0
M1164 363 49 365 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=71300 $D=0
M1165 364 49 366 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=75930 $D=0
M1166 365 361 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=71300 $D=0
M1167 366 362 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=75930 $D=0
M1168 257 367 365 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=71300 $D=0
M1169 258 368 366 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=75930 $D=0
M1170 367 51 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=71300 $D=0
M1171 368 51 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=75930 $D=0
M1172 165 52 369 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=71300 $D=0
M1173 166 52 370 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=75930 $D=0
M1174 371 53 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=71300 $D=0
M1175 372 53 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=75930 $D=0
M1176 373 369 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=71300 $D=0
M1177 374 370 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=75930 $D=0
M1178 165 373 741 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=71300 $D=0
M1179 166 374 742 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=75930 $D=0
M1180 375 741 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=71300 $D=0
M1181 376 742 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=75930 $D=0
M1182 373 52 375 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=71300 $D=0
M1183 374 52 376 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=75930 $D=0
M1184 375 371 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=71300 $D=0
M1185 376 372 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=75930 $D=0
M1186 257 377 375 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=71300 $D=0
M1187 258 378 376 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=75930 $D=0
M1188 377 54 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=71300 $D=0
M1189 378 54 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=75930 $D=0
M1190 165 55 379 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=71300 $D=0
M1191 166 55 380 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=75930 $D=0
M1192 381 56 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=71300 $D=0
M1193 382 56 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=75930 $D=0
M1194 383 379 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=71300 $D=0
M1195 384 380 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=75930 $D=0
M1196 165 383 743 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=71300 $D=0
M1197 166 384 744 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=75930 $D=0
M1198 385 743 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=71300 $D=0
M1199 386 744 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=75930 $D=0
M1200 383 55 385 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=71300 $D=0
M1201 384 55 386 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=75930 $D=0
M1202 385 381 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=71300 $D=0
M1203 386 382 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=75930 $D=0
M1204 257 387 385 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=71300 $D=0
M1205 258 388 386 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=75930 $D=0
M1206 387 57 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=71300 $D=0
M1207 388 57 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=75930 $D=0
M1208 165 58 389 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=71300 $D=0
M1209 166 58 390 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=75930 $D=0
M1210 391 59 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=71300 $D=0
M1211 392 59 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=75930 $D=0
M1212 393 389 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=71300 $D=0
M1213 394 390 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=75930 $D=0
M1214 165 393 745 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=71300 $D=0
M1215 166 394 746 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=75930 $D=0
M1216 395 745 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=71300 $D=0
M1217 396 746 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=75930 $D=0
M1218 393 58 395 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=71300 $D=0
M1219 394 58 396 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=75930 $D=0
M1220 395 391 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=71300 $D=0
M1221 396 392 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=75930 $D=0
M1222 257 397 395 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=71300 $D=0
M1223 258 398 396 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=75930 $D=0
M1224 397 60 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=71300 $D=0
M1225 398 60 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=75930 $D=0
M1226 165 61 399 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=71300 $D=0
M1227 166 61 400 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=75930 $D=0
M1228 401 62 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=71300 $D=0
M1229 402 62 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=75930 $D=0
M1230 403 399 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=71300 $D=0
M1231 404 400 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=75930 $D=0
M1232 165 403 747 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=71300 $D=0
M1233 166 404 748 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=75930 $D=0
M1234 405 747 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=71300 $D=0
M1235 406 748 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=75930 $D=0
M1236 403 61 405 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=71300 $D=0
M1237 404 61 406 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=75930 $D=0
M1238 405 401 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=71300 $D=0
M1239 406 402 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=75930 $D=0
M1240 257 407 405 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=71300 $D=0
M1241 258 408 406 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=75930 $D=0
M1242 407 63 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=71300 $D=0
M1243 408 63 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=75930 $D=0
M1244 165 64 409 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=71300 $D=0
M1245 166 64 410 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=75930 $D=0
M1246 411 65 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=71300 $D=0
M1247 412 65 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=75930 $D=0
M1248 413 409 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=71300 $D=0
M1249 414 410 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=75930 $D=0
M1250 165 413 749 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=71300 $D=0
M1251 166 414 750 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=75930 $D=0
M1252 415 749 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=71300 $D=0
M1253 416 750 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=75930 $D=0
M1254 413 64 415 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=71300 $D=0
M1255 414 64 416 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=75930 $D=0
M1256 415 411 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=71300 $D=0
M1257 416 412 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=75930 $D=0
M1258 257 417 415 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=71300 $D=0
M1259 258 418 416 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=75930 $D=0
M1260 417 66 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=71300 $D=0
M1261 418 66 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=75930 $D=0
M1262 165 67 419 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=71300 $D=0
M1263 166 67 420 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=75930 $D=0
M1264 421 68 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=71300 $D=0
M1265 422 68 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=75930 $D=0
M1266 423 419 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=71300 $D=0
M1267 424 420 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=75930 $D=0
M1268 165 423 751 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=71300 $D=0
M1269 166 424 752 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=75930 $D=0
M1270 425 751 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=71300 $D=0
M1271 426 752 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=75930 $D=0
M1272 423 67 425 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=71300 $D=0
M1273 424 67 426 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=75930 $D=0
M1274 425 421 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=71300 $D=0
M1275 426 422 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=75930 $D=0
M1276 257 427 425 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=71300 $D=0
M1277 258 428 426 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=75930 $D=0
M1278 427 69 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=71300 $D=0
M1279 428 69 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=75930 $D=0
M1280 165 70 429 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=71300 $D=0
M1281 166 70 430 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=75930 $D=0
M1282 431 71 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=71300 $D=0
M1283 432 71 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=75930 $D=0
M1284 433 429 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=71300 $D=0
M1285 434 430 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=75930 $D=0
M1286 165 433 753 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=71300 $D=0
M1287 166 434 754 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=75930 $D=0
M1288 435 753 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=71300 $D=0
M1289 436 754 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=75930 $D=0
M1290 433 70 435 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=71300 $D=0
M1291 434 70 436 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=75930 $D=0
M1292 435 431 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=71300 $D=0
M1293 436 432 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=75930 $D=0
M1294 257 437 435 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=71300 $D=0
M1295 258 438 436 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=75930 $D=0
M1296 437 72 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=71300 $D=0
M1297 438 72 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=75930 $D=0
M1298 165 73 439 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=71300 $D=0
M1299 166 73 440 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=75930 $D=0
M1300 441 74 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=71300 $D=0
M1301 442 74 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=75930 $D=0
M1302 443 439 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=71300 $D=0
M1303 444 440 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=75930 $D=0
M1304 165 443 755 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=71300 $D=0
M1305 166 444 756 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=75930 $D=0
M1306 445 755 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=71300 $D=0
M1307 446 756 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=75930 $D=0
M1308 443 73 445 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=71300 $D=0
M1309 444 73 446 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=75930 $D=0
M1310 445 441 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=71300 $D=0
M1311 446 442 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=75930 $D=0
M1312 257 447 445 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=71300 $D=0
M1313 258 448 446 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=75930 $D=0
M1314 447 75 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=71300 $D=0
M1315 448 75 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=75930 $D=0
M1316 165 76 449 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=71300 $D=0
M1317 166 76 450 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=75930 $D=0
M1318 451 77 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=71300 $D=0
M1319 452 77 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=75930 $D=0
M1320 453 449 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=71300 $D=0
M1321 454 450 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=75930 $D=0
M1322 165 453 757 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=71300 $D=0
M1323 166 454 758 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=75930 $D=0
M1324 455 757 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=71300 $D=0
M1325 456 758 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=75930 $D=0
M1326 453 76 455 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=71300 $D=0
M1327 454 76 456 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=75930 $D=0
M1328 455 451 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=71300 $D=0
M1329 456 452 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=75930 $D=0
M1330 257 457 455 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=71300 $D=0
M1331 258 458 456 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=75930 $D=0
M1332 457 78 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=71300 $D=0
M1333 458 78 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=75930 $D=0
M1334 165 79 459 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=71300 $D=0
M1335 166 79 460 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=75930 $D=0
M1336 461 80 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=71300 $D=0
M1337 462 80 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=75930 $D=0
M1338 463 459 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=71300 $D=0
M1339 464 460 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=75930 $D=0
M1340 165 463 759 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=71300 $D=0
M1341 166 464 760 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=75930 $D=0
M1342 465 759 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=71300 $D=0
M1343 466 760 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=75930 $D=0
M1344 463 79 465 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=71300 $D=0
M1345 464 79 466 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=75930 $D=0
M1346 465 461 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=71300 $D=0
M1347 466 462 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=75930 $D=0
M1348 257 467 465 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=71300 $D=0
M1349 258 468 466 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=75930 $D=0
M1350 467 81 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=71300 $D=0
M1351 468 81 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=75930 $D=0
M1352 165 82 469 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=71300 $D=0
M1353 166 82 470 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=75930 $D=0
M1354 471 83 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=71300 $D=0
M1355 472 83 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=75930 $D=0
M1356 473 469 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=71300 $D=0
M1357 474 470 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=75930 $D=0
M1358 165 473 761 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=71300 $D=0
M1359 166 474 762 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=75930 $D=0
M1360 475 761 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=71300 $D=0
M1361 476 762 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=75930 $D=0
M1362 473 82 475 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=71300 $D=0
M1363 474 82 476 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=75930 $D=0
M1364 475 471 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=71300 $D=0
M1365 476 472 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=75930 $D=0
M1366 257 477 475 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=71300 $D=0
M1367 258 478 476 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=75930 $D=0
M1368 477 84 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=71300 $D=0
M1369 478 84 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=75930 $D=0
M1370 165 85 479 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=71300 $D=0
M1371 166 85 480 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=75930 $D=0
M1372 481 86 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=71300 $D=0
M1373 482 86 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=75930 $D=0
M1374 483 479 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=71300 $D=0
M1375 484 480 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=75930 $D=0
M1376 165 483 763 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=71300 $D=0
M1377 166 484 764 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=75930 $D=0
M1378 485 763 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=71300 $D=0
M1379 486 764 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=75930 $D=0
M1380 483 85 485 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=71300 $D=0
M1381 484 85 486 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=75930 $D=0
M1382 485 481 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=71300 $D=0
M1383 486 482 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=75930 $D=0
M1384 257 487 485 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=71300 $D=0
M1385 258 488 486 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=75930 $D=0
M1386 487 87 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=71300 $D=0
M1387 488 87 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=75930 $D=0
M1388 165 88 489 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=71300 $D=0
M1389 166 88 490 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=75930 $D=0
M1390 491 89 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=71300 $D=0
M1391 492 89 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=75930 $D=0
M1392 493 489 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=71300 $D=0
M1393 494 490 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=75930 $D=0
M1394 165 493 765 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=71300 $D=0
M1395 166 494 766 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=75930 $D=0
M1396 495 765 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=71300 $D=0
M1397 496 766 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=75930 $D=0
M1398 493 88 495 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=71300 $D=0
M1399 494 88 496 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=75930 $D=0
M1400 495 491 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=71300 $D=0
M1401 496 492 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=75930 $D=0
M1402 257 497 495 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=71300 $D=0
M1403 258 498 496 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=75930 $D=0
M1404 497 90 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=71300 $D=0
M1405 498 90 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=75930 $D=0
M1406 165 91 499 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=71300 $D=0
M1407 166 91 500 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=75930 $D=0
M1408 501 92 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=71300 $D=0
M1409 502 92 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=75930 $D=0
M1410 503 499 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=71300 $D=0
M1411 504 500 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=75930 $D=0
M1412 165 503 767 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=71300 $D=0
M1413 166 504 768 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=75930 $D=0
M1414 505 767 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=71300 $D=0
M1415 506 768 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=75930 $D=0
M1416 503 91 505 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=71300 $D=0
M1417 504 91 506 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=75930 $D=0
M1418 505 501 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=71300 $D=0
M1419 506 502 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=75930 $D=0
M1420 257 507 505 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=71300 $D=0
M1421 258 508 506 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=75930 $D=0
M1422 507 93 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=71300 $D=0
M1423 508 93 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=75930 $D=0
M1424 165 94 509 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=71300 $D=0
M1425 166 94 510 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=75930 $D=0
M1426 511 95 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=71300 $D=0
M1427 512 95 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=75930 $D=0
M1428 513 509 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=71300 $D=0
M1429 514 510 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=75930 $D=0
M1430 165 513 769 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=71300 $D=0
M1431 166 514 770 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=75930 $D=0
M1432 515 769 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=71300 $D=0
M1433 516 770 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=75930 $D=0
M1434 513 94 515 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=71300 $D=0
M1435 514 94 516 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=75930 $D=0
M1436 515 511 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=71300 $D=0
M1437 516 512 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=75930 $D=0
M1438 257 517 515 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=71300 $D=0
M1439 258 518 516 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=75930 $D=0
M1440 517 96 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=71300 $D=0
M1441 518 96 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=75930 $D=0
M1442 165 97 519 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=71300 $D=0
M1443 166 97 520 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=75930 $D=0
M1444 521 98 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=71300 $D=0
M1445 522 98 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=75930 $D=0
M1446 523 519 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=71300 $D=0
M1447 524 520 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=75930 $D=0
M1448 165 523 771 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=71300 $D=0
M1449 166 524 772 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=75930 $D=0
M1450 525 771 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=71300 $D=0
M1451 526 772 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=75930 $D=0
M1452 523 97 525 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=71300 $D=0
M1453 524 97 526 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=75930 $D=0
M1454 525 521 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=71300 $D=0
M1455 526 522 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=75930 $D=0
M1456 257 527 525 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=71300 $D=0
M1457 258 528 526 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=75930 $D=0
M1458 527 99 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=71300 $D=0
M1459 528 99 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=75930 $D=0
M1460 165 100 529 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=71300 $D=0
M1461 166 100 530 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=75930 $D=0
M1462 531 101 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=71300 $D=0
M1463 532 101 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=75930 $D=0
M1464 533 529 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=71300 $D=0
M1465 534 530 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=75930 $D=0
M1466 165 533 773 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=71300 $D=0
M1467 166 534 774 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=75930 $D=0
M1468 535 773 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=71300 $D=0
M1469 536 774 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=75930 $D=0
M1470 533 100 535 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=71300 $D=0
M1471 534 100 536 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=75930 $D=0
M1472 535 531 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=71300 $D=0
M1473 536 532 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=75930 $D=0
M1474 257 537 535 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=71300 $D=0
M1475 258 538 536 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=75930 $D=0
M1476 537 102 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=71300 $D=0
M1477 538 102 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=75930 $D=0
M1478 165 103 539 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=71300 $D=0
M1479 166 103 540 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=75930 $D=0
M1480 541 104 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=71300 $D=0
M1481 542 104 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=75930 $D=0
M1482 543 539 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=71300 $D=0
M1483 544 540 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=75930 $D=0
M1484 165 543 775 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=71300 $D=0
M1485 166 544 776 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=75930 $D=0
M1486 545 775 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=71300 $D=0
M1487 546 776 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=75930 $D=0
M1488 543 103 545 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=71300 $D=0
M1489 544 103 546 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=75930 $D=0
M1490 545 541 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=71300 $D=0
M1491 546 542 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=75930 $D=0
M1492 257 547 545 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=71300 $D=0
M1493 258 548 546 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=75930 $D=0
M1494 547 105 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=71300 $D=0
M1495 548 105 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=75930 $D=0
M1496 165 106 549 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=71300 $D=0
M1497 166 106 550 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=75930 $D=0
M1498 551 107 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=71300 $D=0
M1499 552 107 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=75930 $D=0
M1500 553 549 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=71300 $D=0
M1501 554 550 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=75930 $D=0
M1502 165 553 777 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=71300 $D=0
M1503 166 554 778 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=75930 $D=0
M1504 555 777 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=71300 $D=0
M1505 556 778 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=75930 $D=0
M1506 553 106 555 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=71300 $D=0
M1507 554 106 556 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=75930 $D=0
M1508 555 551 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=71300 $D=0
M1509 556 552 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=75930 $D=0
M1510 257 557 555 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=71300 $D=0
M1511 258 558 556 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=75930 $D=0
M1512 557 109 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=71300 $D=0
M1513 558 109 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=75930 $D=0
M1514 165 110 559 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=71300 $D=0
M1515 166 110 560 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=75930 $D=0
M1516 561 111 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=71300 $D=0
M1517 562 111 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=75930 $D=0
M1518 5 561 253 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=71300 $D=0
M1519 6 562 254 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=75930 $D=0
M1520 257 559 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=71300 $D=0
M1521 258 560 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=75930 $D=0
M1522 165 565 563 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=71300 $D=0
M1523 166 566 564 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=75930 $D=0
M1524 565 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=71300 $D=0
M1525 566 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=75930 $D=0
M1526 779 253 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=71300 $D=0
M1527 780 254 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=75930 $D=0
M1528 567 565 779 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=71300 $D=0
M1529 568 566 780 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=75930 $D=0
M1530 165 567 569 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=71300 $D=0
M1531 166 568 570 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=75930 $D=0
M1532 781 569 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=71300 $D=0
M1533 782 570 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=75930 $D=0
M1534 567 563 781 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=71300 $D=0
M1535 568 564 782 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=75930 $D=0
M1536 165 573 571 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=71300 $D=0
M1537 166 574 572 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=75930 $D=0
M1538 573 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=71300 $D=0
M1539 574 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=75930 $D=0
M1540 783 257 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=71300 $D=0
M1541 784 258 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=75930 $D=0
M1542 575 573 783 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=71300 $D=0
M1543 576 574 784 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=75930 $D=0
M1544 165 575 116 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=71300 $D=0
M1545 166 576 117 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=75930 $D=0
M1546 785 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=71300 $D=0
M1547 786 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=75930 $D=0
M1548 575 571 785 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=71300 $D=0
M1549 576 572 786 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=75930 $D=0
M1550 577 120 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=71300 $D=0
M1551 578 120 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=75930 $D=0
M1552 579 120 569 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=71300 $D=0
M1553 580 120 570 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=75930 $D=0
M1554 121 577 579 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=71300 $D=0
M1555 121 578 580 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=75930 $D=0
M1556 581 122 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=71300 $D=0
M1557 582 122 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=75930 $D=0
M1558 583 122 116 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=71300 $D=0
M1559 584 122 117 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=75930 $D=0
M1560 787 581 583 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=71300 $D=0
M1561 788 582 584 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=75930 $D=0
M1562 165 116 787 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=71300 $D=0
M1563 166 117 788 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=75930 $D=0
M1564 585 123 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=71300 $D=0
M1565 586 123 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=75930 $D=0
M1566 587 123 583 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=71300 $D=0
M1567 588 123 584 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=75930 $D=0
M1568 10 585 587 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=71300 $D=0
M1569 11 586 588 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=75930 $D=0
M1570 590 589 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=71300 $D=0
M1571 591 124 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=75930 $D=0
M1572 165 594 592 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=71300 $D=0
M1573 166 595 593 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=75930 $D=0
M1574 596 579 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=71300 $D=0
M1575 597 580 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=75930 $D=0
M1576 594 579 589 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=71300 $D=0
M1577 595 580 124 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=75930 $D=0
M1578 590 596 594 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=71300 $D=0
M1579 591 597 595 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=75930 $D=0
M1580 598 592 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=71300 $D=0
M1581 599 593 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=75930 $D=0
M1582 125 592 587 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=71300 $D=0
M1583 589 593 588 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=75930 $D=0
M1584 579 598 125 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=71300 $D=0
M1585 580 599 589 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=75930 $D=0
M1586 600 125 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=71300 $D=0
M1587 601 589 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=75930 $D=0
M1588 602 592 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=71300 $D=0
M1589 603 593 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=75930 $D=0
M1590 604 592 600 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=71300 $D=0
M1591 605 593 601 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=75930 $D=0
M1592 587 602 604 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=71300 $D=0
M1593 588 603 605 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=75930 $D=0
M1594 799 579 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=70940 $D=0
M1595 800 580 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=75570 $D=0
M1596 606 587 799 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=70940 $D=0
M1597 607 588 800 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=75570 $D=0
M1598 608 604 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=71300 $D=0
M1599 609 605 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=75930 $D=0
M1600 610 579 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=71300 $D=0
M1601 611 580 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=75930 $D=0
M1602 165 587 610 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=71300 $D=0
M1603 166 588 611 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=75930 $D=0
M1604 612 579 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=71300 $D=0
M1605 613 580 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=75930 $D=0
M1606 165 587 612 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=71300 $D=0
M1607 166 588 613 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=75930 $D=0
M1608 801 579 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=71120 $D=0
M1609 802 580 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=75750 $D=0
M1610 616 587 801 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=71120 $D=0
M1611 617 588 802 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=75750 $D=0
M1612 165 612 616 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=71300 $D=0
M1613 166 613 617 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=75930 $D=0
M1614 618 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=71300 $D=0
M1615 619 128 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=75930 $D=0
M1616 620 128 606 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=71300 $D=0
M1617 621 128 607 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=75930 $D=0
M1618 610 618 620 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=71300 $D=0
M1619 611 619 621 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=75930 $D=0
M1620 622 128 608 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=71300 $D=0
M1621 623 128 609 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=75930 $D=0
M1622 616 618 622 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=71300 $D=0
M1623 617 619 623 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=75930 $D=0
M1624 624 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=71300 $D=0
M1625 625 129 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=75930 $D=0
M1626 626 129 622 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=71300 $D=0
M1627 627 129 623 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=75930 $D=0
M1628 620 624 626 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=71300 $D=0
M1629 621 625 627 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=75930 $D=0
M1630 12 626 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=71300 $D=0
M1631 13 627 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=75930 $D=0
M1632 628 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=71300 $D=0
M1633 629 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=75930 $D=0
M1634 630 130 131 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=71300 $D=0
M1635 631 130 132 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=75930 $D=0
M1636 133 628 630 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=71300 $D=0
M1637 134 629 631 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=75930 $D=0
M1638 632 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=71300 $D=0
M1639 633 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=75930 $D=0
M1640 634 130 135 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=71300 $D=0
M1641 635 130 136 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=75930 $D=0
M1642 137 632 634 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=71300 $D=0
M1643 138 633 635 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=75930 $D=0
M1644 636 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=71300 $D=0
M1645 637 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=75930 $D=0
M1646 638 130 126 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=71300 $D=0
M1647 639 130 139 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=75930 $D=0
M1648 114 636 638 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=71300 $D=0
M1649 115 637 639 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=75930 $D=0
M1650 640 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=71300 $D=0
M1651 641 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=75930 $D=0
M1652 642 130 140 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=71300 $D=0
M1653 643 130 141 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=75930 $D=0
M1654 142 640 642 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=71300 $D=0
M1655 143 641 643 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=75930 $D=0
M1656 644 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=71300 $D=0
M1657 645 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=75930 $D=0
M1658 646 130 144 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=71300 $D=0
M1659 647 130 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=75930 $D=0
M1660 145 644 646 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=71300 $D=0
M1661 146 645 647 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=75930 $D=0
M1662 165 579 789 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=71300 $D=0
M1663 166 580 790 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=75930 $D=0
M1664 134 789 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=71300 $D=0
M1665 131 790 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=75930 $D=0
M1666 648 147 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=71300 $D=0
M1667 649 147 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=75930 $D=0
M1668 149 147 134 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=71300 $D=0
M1669 150 147 131 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=75930 $D=0
M1670 630 648 149 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=71300 $D=0
M1671 631 649 150 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=75930 $D=0
M1672 650 151 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=71300 $D=0
M1673 651 151 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=75930 $D=0
M1674 118 151 149 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=71300 $D=0
M1675 119 151 150 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=75930 $D=0
M1676 634 650 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=71300 $D=0
M1677 635 651 119 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=75930 $D=0
M1678 652 152 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=71300 $D=0
M1679 653 152 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=75930 $D=0
M1680 108 152 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=71300 $D=0
M1681 113 152 119 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=75930 $D=0
M1682 638 652 108 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=71300 $D=0
M1683 639 653 113 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=75930 $D=0
M1684 654 153 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=71300 $D=0
M1685 655 153 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=75930 $D=0
M1686 148 153 108 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=71300 $D=0
M1687 154 153 113 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=75930 $D=0
M1688 642 654 148 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=71300 $D=0
M1689 643 655 154 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=75930 $D=0
M1690 656 155 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=71300 $D=0
M1691 657 155 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=75930 $D=0
M1692 229 155 148 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=71300 $D=0
M1693 230 155 154 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=75930 $D=0
M1694 646 656 229 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=71300 $D=0
M1695 647 657 230 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=75930 $D=0
M1696 658 156 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=71300 $D=0
M1697 659 156 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=75930 $D=0
M1698 660 156 116 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=71300 $D=0
M1699 661 156 117 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=75930 $D=0
M1700 10 658 660 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=71300 $D=0
M1701 11 659 661 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=75930 $D=0
M1702 662 569 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=71300 $D=0
M1703 663 570 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=75930 $D=0
M1704 165 660 662 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=71300 $D=0
M1705 166 661 663 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=75930 $D=0
M1706 803 569 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=71120 $D=0
M1707 804 570 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=75750 $D=0
M1708 666 660 803 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=71120 $D=0
M1709 667 661 804 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=75750 $D=0
M1710 165 662 666 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=71300 $D=0
M1711 166 663 667 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=75930 $D=0
M1712 791 157 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=71300 $D=0
M1713 792 668 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=75930 $D=0
M1714 165 666 791 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=71300 $D=0
M1715 166 667 792 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=75930 $D=0
M1716 668 791 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=71300 $D=0
M1717 158 792 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=75930 $D=0
M1718 805 569 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=70940 $D=0
M1719 806 570 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=75570 $D=0
M1720 669 671 805 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=70940 $D=0
M1721 670 672 806 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=75570 $D=0
M1722 671 660 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=71300 $D=0
M1723 672 661 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=75930 $D=0
M1724 673 669 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=71300 $D=0
M1725 674 670 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=75930 $D=0
M1726 165 157 673 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=71300 $D=0
M1727 166 668 674 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=75930 $D=0
M1728 676 159 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=71300 $D=0
M1729 677 675 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=75930 $D=0
M1730 675 673 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=71300 $D=0
M1731 160 674 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=75930 $D=0
M1732 165 676 675 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=71300 $D=0
M1733 166 677 160 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=75930 $D=0
M1734 679 678 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=71300 $D=0
M1735 680 161 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=75930 $D=0
M1736 165 683 681 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=71300 $D=0
M1737 166 684 682 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=75930 $D=0
M1738 685 121 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=71300 $D=0
M1739 686 121 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=75930 $D=0
M1740 683 121 678 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=71300 $D=0
M1741 684 121 161 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=75930 $D=0
M1742 679 685 683 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=71300 $D=0
M1743 680 686 684 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=75930 $D=0
M1744 687 681 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=71300 $D=0
M1745 688 682 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=75930 $D=0
M1746 162 681 5 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=71300 $D=0
M1747 678 682 6 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=75930 $D=0
M1748 121 687 162 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=71300 $D=0
M1749 121 688 678 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=75930 $D=0
M1750 689 162 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=71300 $D=0
M1751 690 678 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=75930 $D=0
M1752 691 681 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=71300 $D=0
M1753 692 682 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=75930 $D=0
M1754 231 681 689 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=71300 $D=0
M1755 232 682 690 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=75930 $D=0
M1756 5 691 231 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=71300 $D=0
M1757 6 692 232 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=75930 $D=0
M1758 693 163 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=71300 $D=0
M1759 694 163 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=75930 $D=0
M1760 695 163 231 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=71300 $D=0
M1761 696 163 232 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=75930 $D=0
M1762 12 693 695 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=71300 $D=0
M1763 13 694 696 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=75930 $D=0
M1764 697 164 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=71300 $D=0
M1765 698 164 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=75930 $D=0
M1766 164 164 695 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=71300 $D=0
M1767 164 164 696 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=75930 $D=0
M1768 5 697 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=71300 $D=0
M1769 6 698 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=75930 $D=0
M1770 699 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=71300 $D=0
M1771 700 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=75930 $D=0
M1772 165 699 701 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=71300 $D=0
M1773 166 700 702 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=75930 $D=0
M1774 703 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=71300 $D=0
M1775 704 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=75930 $D=0
M1776 705 701 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=71300 $D=0
M1777 706 702 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=75930 $D=0
M1778 165 705 793 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=71300 $D=0
M1779 166 706 794 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=75930 $D=0
M1780 707 793 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=71300 $D=0
M1781 708 794 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=75930 $D=0
M1782 705 699 707 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=71300 $D=0
M1783 706 700 708 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=75930 $D=0
M1784 709 703 707 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=71300 $D=0
M1785 710 704 708 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=75930 $D=0
M1786 165 713 711 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=71300 $D=0
M1787 166 714 712 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=75930 $D=0
M1788 713 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=71300 $D=0
M1789 714 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=75930 $D=0
M1790 795 709 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=71300 $D=0
M1791 796 710 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=75930 $D=0
M1792 715 713 795 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=71300 $D=0
M1793 716 714 796 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=75930 $D=0
M1794 165 715 121 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=71300 $D=0
M1795 166 716 121 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=75930 $D=0
M1796 797 121 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=71300 $D=0
M1797 798 121 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=75930 $D=0
M1798 715 711 797 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=71300 $D=0
M1799 716 712 798 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=75930 $D=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194
** N=1452 EP=194 IP=2964 FDC=3600
M0 221 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=51530 $D=1
M1 222 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=56160 $D=1
M2 223 1 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=60790 $D=1
M3 224 1 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=65420 $D=1
M4 225 221 2 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=51530 $D=1
M5 226 222 3 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=56160 $D=1
M6 227 223 4 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=60790 $D=1
M7 228 224 5 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=65420 $D=1
M8 8 1 225 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=51530 $D=1
M9 9 1 226 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=56160 $D=1
M10 10 1 227 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=60790 $D=1
M11 11 1 228 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=65420 $D=1
M12 229 221 6 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=51530 $D=1
M13 230 222 6 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=56160 $D=1
M14 231 223 6 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=60790 $D=1
M15 232 224 6 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=65420 $D=1
M16 7 1 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=51530 $D=1
M17 7 1 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=56160 $D=1
M18 7 1 231 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=60790 $D=1
M19 7 1 232 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=65420 $D=1
M20 233 221 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=51530 $D=1
M21 234 222 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=56160 $D=1
M22 235 223 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=60790 $D=1
M23 236 224 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=65420 $D=1
M24 8 1 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=51530 $D=1
M25 9 1 234 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=56160 $D=1
M26 10 1 235 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=60790 $D=1
M27 11 1 236 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=65420 $D=1
M28 241 237 233 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=51530 $D=1
M29 242 238 234 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=56160 $D=1
M30 243 239 235 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=60790 $D=1
M31 244 240 236 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=65420 $D=1
M32 237 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=51530 $D=1
M33 238 12 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=56160 $D=1
M34 239 12 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=60790 $D=1
M35 240 12 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=65420 $D=1
M36 245 237 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=51530 $D=1
M37 246 238 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=56160 $D=1
M38 247 239 231 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=60790 $D=1
M39 248 240 232 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=65420 $D=1
M40 225 12 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=51530 $D=1
M41 226 12 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=56160 $D=1
M42 227 12 247 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=60790 $D=1
M43 228 12 248 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=65420 $D=1
M44 249 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=51530 $D=1
M45 250 13 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=56160 $D=1
M46 251 13 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=60790 $D=1
M47 252 13 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=65420 $D=1
M48 253 249 245 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=51530 $D=1
M49 254 250 246 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=56160 $D=1
M50 255 251 247 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=60790 $D=1
M51 256 252 248 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=65420 $D=1
M52 241 13 253 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=51530 $D=1
M53 242 13 254 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=56160 $D=1
M54 243 13 255 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=60790 $D=1
M55 244 13 256 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=65420 $D=1
M56 257 14 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=51530 $D=1
M57 258 14 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=56160 $D=1
M58 259 14 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=60790 $D=1
M59 260 14 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=65420 $D=1
M60 261 257 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=51530 $D=1
M61 262 258 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=56160 $D=1
M62 263 259 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=60790 $D=1
M63 264 260 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=65420 $D=1
M64 15 14 261 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=51530 $D=1
M65 16 14 262 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=56160 $D=1
M66 17 14 263 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=60790 $D=1
M67 18 14 264 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=65420 $D=1
M68 265 257 19 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=51530 $D=1
M69 266 258 20 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=56160 $D=1
M70 267 259 21 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=60790 $D=1
M71 268 260 22 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=65420 $D=1
M72 269 14 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=51530 $D=1
M73 270 14 266 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=56160 $D=1
M74 271 14 267 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=60790 $D=1
M75 272 14 268 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=65420 $D=1
M76 277 257 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=51530 $D=1
M77 278 258 274 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=56160 $D=1
M78 279 259 275 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=60790 $D=1
M79 280 260 276 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=65420 $D=1
M80 253 14 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=51530 $D=1
M81 254 14 278 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=56160 $D=1
M82 255 14 279 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=60790 $D=1
M83 256 14 280 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=65420 $D=1
M84 285 281 277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=51530 $D=1
M85 286 282 278 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=56160 $D=1
M86 287 283 279 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=60790 $D=1
M87 288 284 280 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=65420 $D=1
M88 281 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=51530 $D=1
M89 282 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=56160 $D=1
M90 283 23 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=60790 $D=1
M91 284 23 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=65420 $D=1
M92 289 281 265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=51530 $D=1
M93 290 282 266 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=56160 $D=1
M94 291 283 267 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=60790 $D=1
M95 292 284 268 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=65420 $D=1
M96 261 23 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=51530 $D=1
M97 262 23 290 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=56160 $D=1
M98 263 23 291 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=60790 $D=1
M99 264 23 292 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=65420 $D=1
M100 293 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=51530 $D=1
M101 294 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=56160 $D=1
M102 295 24 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=60790 $D=1
M103 296 24 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=65420 $D=1
M104 297 293 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=51530 $D=1
M105 298 294 290 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=56160 $D=1
M106 299 295 291 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=60790 $D=1
M107 300 296 292 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=65420 $D=1
M108 285 24 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=51530 $D=1
M109 286 24 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=56160 $D=1
M110 287 24 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=60790 $D=1
M111 288 24 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=65420 $D=1
M112 8 25 301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=51530 $D=1
M113 9 25 302 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=56160 $D=1
M114 10 25 303 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=60790 $D=1
M115 11 25 304 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=65420 $D=1
M116 305 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=51530 $D=1
M117 306 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=56160 $D=1
M118 307 26 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=60790 $D=1
M119 308 26 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=65420 $D=1
M120 309 25 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=51530 $D=1
M121 310 25 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=56160 $D=1
M122 311 25 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=60790 $D=1
M123 312 25 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=65420 $D=1
M124 8 309 1249 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=51530 $D=1
M125 9 310 1250 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=56160 $D=1
M126 10 311 1251 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=60790 $D=1
M127 11 312 1252 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=65420 $D=1
M128 313 1249 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=51530 $D=1
M129 314 1250 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=56160 $D=1
M130 315 1251 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=60790 $D=1
M131 316 1252 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=65420 $D=1
M132 309 301 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=51530 $D=1
M133 310 302 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=56160 $D=1
M134 311 303 315 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=60790 $D=1
M135 312 304 316 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=65420 $D=1
M136 313 26 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=51530 $D=1
M137 314 26 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=56160 $D=1
M138 315 26 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=60790 $D=1
M139 316 26 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=65420 $D=1
M140 325 27 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=51530 $D=1
M141 326 27 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=56160 $D=1
M142 327 27 315 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=60790 $D=1
M143 328 27 316 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=65420 $D=1
M144 321 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=51530 $D=1
M145 322 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=56160 $D=1
M146 323 27 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=60790 $D=1
M147 324 27 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=65420 $D=1
M148 8 28 329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=51530 $D=1
M149 9 28 330 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=56160 $D=1
M150 10 28 331 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=60790 $D=1
M151 11 28 332 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=65420 $D=1
M152 333 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=51530 $D=1
M153 334 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=56160 $D=1
M154 335 29 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=60790 $D=1
M155 336 29 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=65420 $D=1
M156 337 28 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=51530 $D=1
M157 338 28 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=56160 $D=1
M158 339 28 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=60790 $D=1
M159 340 28 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=65420 $D=1
M160 8 337 1253 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=51530 $D=1
M161 9 338 1254 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=56160 $D=1
M162 10 339 1255 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=60790 $D=1
M163 11 340 1256 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=65420 $D=1
M164 341 1253 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=51530 $D=1
M165 342 1254 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=56160 $D=1
M166 343 1255 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=60790 $D=1
M167 344 1256 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=65420 $D=1
M168 337 329 341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=51530 $D=1
M169 338 330 342 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=56160 $D=1
M170 339 331 343 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=60790 $D=1
M171 340 332 344 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=65420 $D=1
M172 341 29 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=51530 $D=1
M173 342 29 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=56160 $D=1
M174 343 29 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=60790 $D=1
M175 344 29 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=65420 $D=1
M176 325 30 341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=51530 $D=1
M177 326 30 342 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=56160 $D=1
M178 327 30 343 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=60790 $D=1
M179 328 30 344 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=65420 $D=1
M180 345 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=51530 $D=1
M181 346 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=56160 $D=1
M182 347 30 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=60790 $D=1
M183 348 30 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=65420 $D=1
M184 8 31 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=51530 $D=1
M185 9 31 350 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=56160 $D=1
M186 10 31 351 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=60790 $D=1
M187 11 31 352 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=65420 $D=1
M188 353 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=51530 $D=1
M189 354 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=56160 $D=1
M190 355 32 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=60790 $D=1
M191 356 32 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=65420 $D=1
M192 357 31 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=51530 $D=1
M193 358 31 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=56160 $D=1
M194 359 31 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=60790 $D=1
M195 360 31 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=65420 $D=1
M196 8 357 1257 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=51530 $D=1
M197 9 358 1258 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=56160 $D=1
M198 10 359 1259 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=60790 $D=1
M199 11 360 1260 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=65420 $D=1
M200 361 1257 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=51530 $D=1
M201 362 1258 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=56160 $D=1
M202 363 1259 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=60790 $D=1
M203 364 1260 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=65420 $D=1
M204 357 349 361 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=51530 $D=1
M205 358 350 362 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=56160 $D=1
M206 359 351 363 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=60790 $D=1
M207 360 352 364 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=65420 $D=1
M208 361 32 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=51530 $D=1
M209 362 32 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=56160 $D=1
M210 363 32 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=60790 $D=1
M211 364 32 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=65420 $D=1
M212 325 33 361 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=51530 $D=1
M213 326 33 362 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=56160 $D=1
M214 327 33 363 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=60790 $D=1
M215 328 33 364 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=65420 $D=1
M216 365 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=51530 $D=1
M217 366 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=56160 $D=1
M218 367 33 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=60790 $D=1
M219 368 33 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=65420 $D=1
M220 8 34 369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=51530 $D=1
M221 9 34 370 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=56160 $D=1
M222 10 34 371 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=60790 $D=1
M223 11 34 372 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=65420 $D=1
M224 373 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=51530 $D=1
M225 374 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=56160 $D=1
M226 375 35 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=60790 $D=1
M227 376 35 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=65420 $D=1
M228 377 34 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=51530 $D=1
M229 378 34 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=56160 $D=1
M230 379 34 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=60790 $D=1
M231 380 34 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=65420 $D=1
M232 8 377 1261 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=51530 $D=1
M233 9 378 1262 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=56160 $D=1
M234 10 379 1263 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=60790 $D=1
M235 11 380 1264 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=65420 $D=1
M236 381 1261 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=51530 $D=1
M237 382 1262 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=56160 $D=1
M238 383 1263 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=60790 $D=1
M239 384 1264 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=65420 $D=1
M240 377 369 381 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=51530 $D=1
M241 378 370 382 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=56160 $D=1
M242 379 371 383 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=60790 $D=1
M243 380 372 384 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=65420 $D=1
M244 381 35 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=51530 $D=1
M245 382 35 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=56160 $D=1
M246 383 35 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=60790 $D=1
M247 384 35 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=65420 $D=1
M248 325 36 381 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=51530 $D=1
M249 326 36 382 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=56160 $D=1
M250 327 36 383 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=60790 $D=1
M251 328 36 384 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=65420 $D=1
M252 385 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=51530 $D=1
M253 386 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=56160 $D=1
M254 387 36 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=60790 $D=1
M255 388 36 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=65420 $D=1
M256 8 37 389 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=51530 $D=1
M257 9 37 390 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=56160 $D=1
M258 10 37 391 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=60790 $D=1
M259 11 37 392 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=65420 $D=1
M260 393 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=51530 $D=1
M261 394 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=56160 $D=1
M262 395 38 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=60790 $D=1
M263 396 38 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=65420 $D=1
M264 397 37 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=51530 $D=1
M265 398 37 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=56160 $D=1
M266 399 37 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=60790 $D=1
M267 400 37 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=65420 $D=1
M268 8 397 1265 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=51530 $D=1
M269 9 398 1266 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=56160 $D=1
M270 10 399 1267 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=60790 $D=1
M271 11 400 1268 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=65420 $D=1
M272 401 1265 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=51530 $D=1
M273 402 1266 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=56160 $D=1
M274 403 1267 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=60790 $D=1
M275 404 1268 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=65420 $D=1
M276 397 389 401 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=51530 $D=1
M277 398 390 402 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=56160 $D=1
M278 399 391 403 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=60790 $D=1
M279 400 392 404 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=65420 $D=1
M280 401 38 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=51530 $D=1
M281 402 38 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=56160 $D=1
M282 403 38 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=60790 $D=1
M283 404 38 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=65420 $D=1
M284 325 39 401 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=51530 $D=1
M285 326 39 402 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=56160 $D=1
M286 327 39 403 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=60790 $D=1
M287 328 39 404 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=65420 $D=1
M288 405 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=51530 $D=1
M289 406 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=56160 $D=1
M290 407 39 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=60790 $D=1
M291 408 39 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=65420 $D=1
M292 8 40 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=51530 $D=1
M293 9 40 410 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=56160 $D=1
M294 10 40 411 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=60790 $D=1
M295 11 40 412 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=65420 $D=1
M296 413 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=51530 $D=1
M297 414 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=56160 $D=1
M298 415 41 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=60790 $D=1
M299 416 41 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=65420 $D=1
M300 417 40 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=51530 $D=1
M301 418 40 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=56160 $D=1
M302 419 40 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=60790 $D=1
M303 420 40 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=65420 $D=1
M304 8 417 1269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=51530 $D=1
M305 9 418 1270 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=56160 $D=1
M306 10 419 1271 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=60790 $D=1
M307 11 420 1272 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=65420 $D=1
M308 421 1269 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=51530 $D=1
M309 422 1270 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=56160 $D=1
M310 423 1271 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=60790 $D=1
M311 424 1272 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=65420 $D=1
M312 417 409 421 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=51530 $D=1
M313 418 410 422 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=56160 $D=1
M314 419 411 423 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=60790 $D=1
M315 420 412 424 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=65420 $D=1
M316 421 41 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=51530 $D=1
M317 422 41 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=56160 $D=1
M318 423 41 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=60790 $D=1
M319 424 41 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=65420 $D=1
M320 325 42 421 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=51530 $D=1
M321 326 42 422 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=56160 $D=1
M322 327 42 423 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=60790 $D=1
M323 328 42 424 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=65420 $D=1
M324 425 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=51530 $D=1
M325 426 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=56160 $D=1
M326 427 42 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=60790 $D=1
M327 428 42 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=65420 $D=1
M328 8 43 429 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=51530 $D=1
M329 9 43 430 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=56160 $D=1
M330 10 43 431 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=60790 $D=1
M331 11 43 432 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=65420 $D=1
M332 433 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=51530 $D=1
M333 434 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=56160 $D=1
M334 435 44 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=60790 $D=1
M335 436 44 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=65420 $D=1
M336 437 43 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=51530 $D=1
M337 438 43 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=56160 $D=1
M338 439 43 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=60790 $D=1
M339 440 43 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=65420 $D=1
M340 8 437 1273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=51530 $D=1
M341 9 438 1274 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=56160 $D=1
M342 10 439 1275 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=60790 $D=1
M343 11 440 1276 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=65420 $D=1
M344 441 1273 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=51530 $D=1
M345 442 1274 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=56160 $D=1
M346 443 1275 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=60790 $D=1
M347 444 1276 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=65420 $D=1
M348 437 429 441 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=51530 $D=1
M349 438 430 442 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=56160 $D=1
M350 439 431 443 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=60790 $D=1
M351 440 432 444 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=65420 $D=1
M352 441 44 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=51530 $D=1
M353 442 44 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=56160 $D=1
M354 443 44 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=60790 $D=1
M355 444 44 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=65420 $D=1
M356 325 45 441 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=51530 $D=1
M357 326 45 442 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=56160 $D=1
M358 327 45 443 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=60790 $D=1
M359 328 45 444 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=65420 $D=1
M360 445 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=51530 $D=1
M361 446 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=56160 $D=1
M362 447 45 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=60790 $D=1
M363 448 45 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=65420 $D=1
M364 8 46 449 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=51530 $D=1
M365 9 46 450 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=56160 $D=1
M366 10 46 451 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=60790 $D=1
M367 11 46 452 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=65420 $D=1
M368 453 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=51530 $D=1
M369 454 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=56160 $D=1
M370 455 47 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=60790 $D=1
M371 456 47 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=65420 $D=1
M372 457 46 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=51530 $D=1
M373 458 46 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=56160 $D=1
M374 459 46 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=60790 $D=1
M375 460 46 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=65420 $D=1
M376 8 457 1277 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=51530 $D=1
M377 9 458 1278 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=56160 $D=1
M378 10 459 1279 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=60790 $D=1
M379 11 460 1280 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=65420 $D=1
M380 461 1277 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=51530 $D=1
M381 462 1278 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=56160 $D=1
M382 463 1279 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=60790 $D=1
M383 464 1280 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=65420 $D=1
M384 457 449 461 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=51530 $D=1
M385 458 450 462 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=56160 $D=1
M386 459 451 463 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=60790 $D=1
M387 460 452 464 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=65420 $D=1
M388 461 47 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=51530 $D=1
M389 462 47 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=56160 $D=1
M390 463 47 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=60790 $D=1
M391 464 47 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=65420 $D=1
M392 325 48 461 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=51530 $D=1
M393 326 48 462 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=56160 $D=1
M394 327 48 463 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=60790 $D=1
M395 328 48 464 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=65420 $D=1
M396 465 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=51530 $D=1
M397 466 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=56160 $D=1
M398 467 48 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=60790 $D=1
M399 468 48 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=65420 $D=1
M400 8 49 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=51530 $D=1
M401 9 49 470 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=56160 $D=1
M402 10 49 471 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=60790 $D=1
M403 11 49 472 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=65420 $D=1
M404 473 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=51530 $D=1
M405 474 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=56160 $D=1
M406 475 50 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=60790 $D=1
M407 476 50 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=65420 $D=1
M408 477 49 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=51530 $D=1
M409 478 49 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=56160 $D=1
M410 479 49 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=60790 $D=1
M411 480 49 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=65420 $D=1
M412 8 477 1281 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=51530 $D=1
M413 9 478 1282 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=56160 $D=1
M414 10 479 1283 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=60790 $D=1
M415 11 480 1284 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=65420 $D=1
M416 481 1281 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=51530 $D=1
M417 482 1282 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=56160 $D=1
M418 483 1283 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=60790 $D=1
M419 484 1284 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=65420 $D=1
M420 477 469 481 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=51530 $D=1
M421 478 470 482 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=56160 $D=1
M422 479 471 483 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=60790 $D=1
M423 480 472 484 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=65420 $D=1
M424 481 50 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=51530 $D=1
M425 482 50 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=56160 $D=1
M426 483 50 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=60790 $D=1
M427 484 50 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=65420 $D=1
M428 325 51 481 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=51530 $D=1
M429 326 51 482 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=56160 $D=1
M430 327 51 483 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=60790 $D=1
M431 328 51 484 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=65420 $D=1
M432 485 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=51530 $D=1
M433 486 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=56160 $D=1
M434 487 51 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=60790 $D=1
M435 488 51 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=65420 $D=1
M436 8 52 489 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=51530 $D=1
M437 9 52 490 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=56160 $D=1
M438 10 52 491 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=60790 $D=1
M439 11 52 492 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=65420 $D=1
M440 493 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=51530 $D=1
M441 494 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=56160 $D=1
M442 495 53 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=60790 $D=1
M443 496 53 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=65420 $D=1
M444 497 52 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=51530 $D=1
M445 498 52 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=56160 $D=1
M446 499 52 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=60790 $D=1
M447 500 52 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=65420 $D=1
M448 8 497 1285 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=51530 $D=1
M449 9 498 1286 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=56160 $D=1
M450 10 499 1287 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=60790 $D=1
M451 11 500 1288 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=65420 $D=1
M452 501 1285 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=51530 $D=1
M453 502 1286 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=56160 $D=1
M454 503 1287 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=60790 $D=1
M455 504 1288 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=65420 $D=1
M456 497 489 501 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=51530 $D=1
M457 498 490 502 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=56160 $D=1
M458 499 491 503 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=60790 $D=1
M459 500 492 504 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=65420 $D=1
M460 501 53 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=51530 $D=1
M461 502 53 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=56160 $D=1
M462 503 53 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=60790 $D=1
M463 504 53 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=65420 $D=1
M464 325 54 501 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=51530 $D=1
M465 326 54 502 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=56160 $D=1
M466 327 54 503 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=60790 $D=1
M467 328 54 504 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=65420 $D=1
M468 505 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=51530 $D=1
M469 506 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=56160 $D=1
M470 507 54 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=60790 $D=1
M471 508 54 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=65420 $D=1
M472 8 55 509 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=51530 $D=1
M473 9 55 510 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=56160 $D=1
M474 10 55 511 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=60790 $D=1
M475 11 55 512 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=65420 $D=1
M476 513 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=51530 $D=1
M477 514 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=56160 $D=1
M478 515 56 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=60790 $D=1
M479 516 56 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=65420 $D=1
M480 517 55 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=51530 $D=1
M481 518 55 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=56160 $D=1
M482 519 55 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=60790 $D=1
M483 520 55 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=65420 $D=1
M484 8 517 1289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=51530 $D=1
M485 9 518 1290 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=56160 $D=1
M486 10 519 1291 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=60790 $D=1
M487 11 520 1292 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=65420 $D=1
M488 521 1289 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=51530 $D=1
M489 522 1290 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=56160 $D=1
M490 523 1291 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=60790 $D=1
M491 524 1292 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=65420 $D=1
M492 517 509 521 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=51530 $D=1
M493 518 510 522 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=56160 $D=1
M494 519 511 523 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=60790 $D=1
M495 520 512 524 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=65420 $D=1
M496 521 56 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=51530 $D=1
M497 522 56 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=56160 $D=1
M498 523 56 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=60790 $D=1
M499 524 56 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=65420 $D=1
M500 325 57 521 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=51530 $D=1
M501 326 57 522 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=56160 $D=1
M502 327 57 523 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=60790 $D=1
M503 328 57 524 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=65420 $D=1
M504 525 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=51530 $D=1
M505 526 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=56160 $D=1
M506 527 57 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=60790 $D=1
M507 528 57 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=65420 $D=1
M508 8 58 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=51530 $D=1
M509 9 58 530 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=56160 $D=1
M510 10 58 531 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=60790 $D=1
M511 11 58 532 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=65420 $D=1
M512 533 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=51530 $D=1
M513 534 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=56160 $D=1
M514 535 59 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=60790 $D=1
M515 536 59 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=65420 $D=1
M516 537 58 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=51530 $D=1
M517 538 58 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=56160 $D=1
M518 539 58 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=60790 $D=1
M519 540 58 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=65420 $D=1
M520 8 537 1293 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=51530 $D=1
M521 9 538 1294 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=56160 $D=1
M522 10 539 1295 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=60790 $D=1
M523 11 540 1296 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=65420 $D=1
M524 541 1293 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=51530 $D=1
M525 542 1294 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=56160 $D=1
M526 543 1295 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=60790 $D=1
M527 544 1296 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=65420 $D=1
M528 537 529 541 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=51530 $D=1
M529 538 530 542 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=56160 $D=1
M530 539 531 543 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=60790 $D=1
M531 540 532 544 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=65420 $D=1
M532 541 59 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=51530 $D=1
M533 542 59 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=56160 $D=1
M534 543 59 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=60790 $D=1
M535 544 59 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=65420 $D=1
M536 325 60 541 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=51530 $D=1
M537 326 60 542 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=56160 $D=1
M538 327 60 543 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=60790 $D=1
M539 328 60 544 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=65420 $D=1
M540 545 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=51530 $D=1
M541 546 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=56160 $D=1
M542 547 60 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=60790 $D=1
M543 548 60 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=65420 $D=1
M544 8 61 549 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=51530 $D=1
M545 9 61 550 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=56160 $D=1
M546 10 61 551 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=60790 $D=1
M547 11 61 552 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=65420 $D=1
M548 553 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=51530 $D=1
M549 554 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=56160 $D=1
M550 555 62 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=60790 $D=1
M551 556 62 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=65420 $D=1
M552 557 61 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=51530 $D=1
M553 558 61 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=56160 $D=1
M554 559 61 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=60790 $D=1
M555 560 61 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=65420 $D=1
M556 8 557 1297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=51530 $D=1
M557 9 558 1298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=56160 $D=1
M558 10 559 1299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=60790 $D=1
M559 11 560 1300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=65420 $D=1
M560 561 1297 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=51530 $D=1
M561 562 1298 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=56160 $D=1
M562 563 1299 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=60790 $D=1
M563 564 1300 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=65420 $D=1
M564 557 549 561 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=51530 $D=1
M565 558 550 562 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=56160 $D=1
M566 559 551 563 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=60790 $D=1
M567 560 552 564 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=65420 $D=1
M568 561 62 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=51530 $D=1
M569 562 62 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=56160 $D=1
M570 563 62 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=60790 $D=1
M571 564 62 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=65420 $D=1
M572 325 63 561 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=51530 $D=1
M573 326 63 562 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=56160 $D=1
M574 327 63 563 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=60790 $D=1
M575 328 63 564 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=65420 $D=1
M576 565 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=51530 $D=1
M577 566 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=56160 $D=1
M578 567 63 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=60790 $D=1
M579 568 63 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=65420 $D=1
M580 8 64 569 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=51530 $D=1
M581 9 64 570 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=56160 $D=1
M582 10 64 571 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=60790 $D=1
M583 11 64 572 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=65420 $D=1
M584 573 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=51530 $D=1
M585 574 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=56160 $D=1
M586 575 65 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=60790 $D=1
M587 576 65 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=65420 $D=1
M588 577 64 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=51530 $D=1
M589 578 64 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=56160 $D=1
M590 579 64 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=60790 $D=1
M591 580 64 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=65420 $D=1
M592 8 577 1301 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=51530 $D=1
M593 9 578 1302 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=56160 $D=1
M594 10 579 1303 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=60790 $D=1
M595 11 580 1304 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=65420 $D=1
M596 581 1301 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=51530 $D=1
M597 582 1302 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=56160 $D=1
M598 583 1303 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=60790 $D=1
M599 584 1304 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=65420 $D=1
M600 577 569 581 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=51530 $D=1
M601 578 570 582 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=56160 $D=1
M602 579 571 583 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=60790 $D=1
M603 580 572 584 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=65420 $D=1
M604 581 65 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=51530 $D=1
M605 582 65 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=56160 $D=1
M606 583 65 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=60790 $D=1
M607 584 65 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=65420 $D=1
M608 325 66 581 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=51530 $D=1
M609 326 66 582 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=56160 $D=1
M610 327 66 583 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=60790 $D=1
M611 328 66 584 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=65420 $D=1
M612 585 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=51530 $D=1
M613 586 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=56160 $D=1
M614 587 66 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=60790 $D=1
M615 588 66 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=65420 $D=1
M616 8 67 589 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=51530 $D=1
M617 9 67 590 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=56160 $D=1
M618 10 67 591 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=60790 $D=1
M619 11 67 592 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=65420 $D=1
M620 593 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=51530 $D=1
M621 594 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=56160 $D=1
M622 595 68 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=60790 $D=1
M623 596 68 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=65420 $D=1
M624 597 67 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=51530 $D=1
M625 598 67 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=56160 $D=1
M626 599 67 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=60790 $D=1
M627 600 67 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=65420 $D=1
M628 8 597 1305 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=51530 $D=1
M629 9 598 1306 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=56160 $D=1
M630 10 599 1307 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=60790 $D=1
M631 11 600 1308 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=65420 $D=1
M632 601 1305 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=51530 $D=1
M633 602 1306 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=56160 $D=1
M634 603 1307 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=60790 $D=1
M635 604 1308 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=65420 $D=1
M636 597 589 601 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=51530 $D=1
M637 598 590 602 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=56160 $D=1
M638 599 591 603 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=60790 $D=1
M639 600 592 604 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=65420 $D=1
M640 601 68 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=51530 $D=1
M641 602 68 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=56160 $D=1
M642 603 68 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=60790 $D=1
M643 604 68 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=65420 $D=1
M644 325 69 601 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=51530 $D=1
M645 326 69 602 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=56160 $D=1
M646 327 69 603 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=60790 $D=1
M647 328 69 604 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=65420 $D=1
M648 605 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=51530 $D=1
M649 606 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=56160 $D=1
M650 607 69 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=60790 $D=1
M651 608 69 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=65420 $D=1
M652 8 70 609 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=51530 $D=1
M653 9 70 610 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=56160 $D=1
M654 10 70 611 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=60790 $D=1
M655 11 70 612 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=65420 $D=1
M656 613 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=51530 $D=1
M657 614 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=56160 $D=1
M658 615 71 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=60790 $D=1
M659 616 71 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=65420 $D=1
M660 617 70 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=51530 $D=1
M661 618 70 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=56160 $D=1
M662 619 70 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=60790 $D=1
M663 620 70 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=65420 $D=1
M664 8 617 1309 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=51530 $D=1
M665 9 618 1310 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=56160 $D=1
M666 10 619 1311 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=60790 $D=1
M667 11 620 1312 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=65420 $D=1
M668 621 1309 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=51530 $D=1
M669 622 1310 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=56160 $D=1
M670 623 1311 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=60790 $D=1
M671 624 1312 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=65420 $D=1
M672 617 609 621 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=51530 $D=1
M673 618 610 622 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=56160 $D=1
M674 619 611 623 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=60790 $D=1
M675 620 612 624 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=65420 $D=1
M676 621 71 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=51530 $D=1
M677 622 71 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=56160 $D=1
M678 623 71 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=60790 $D=1
M679 624 71 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=65420 $D=1
M680 325 72 621 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=51530 $D=1
M681 326 72 622 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=56160 $D=1
M682 327 72 623 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=60790 $D=1
M683 328 72 624 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=65420 $D=1
M684 625 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=51530 $D=1
M685 626 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=56160 $D=1
M686 627 72 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=60790 $D=1
M687 628 72 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=65420 $D=1
M688 8 73 629 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=51530 $D=1
M689 9 73 630 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=56160 $D=1
M690 10 73 631 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=60790 $D=1
M691 11 73 632 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=65420 $D=1
M692 633 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=51530 $D=1
M693 634 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=56160 $D=1
M694 635 74 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=60790 $D=1
M695 636 74 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=65420 $D=1
M696 637 73 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=51530 $D=1
M697 638 73 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=56160 $D=1
M698 639 73 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=60790 $D=1
M699 640 73 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=65420 $D=1
M700 8 637 1313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=51530 $D=1
M701 9 638 1314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=56160 $D=1
M702 10 639 1315 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=60790 $D=1
M703 11 640 1316 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=65420 $D=1
M704 641 1313 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=51530 $D=1
M705 642 1314 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=56160 $D=1
M706 643 1315 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=60790 $D=1
M707 644 1316 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=65420 $D=1
M708 637 629 641 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=51530 $D=1
M709 638 630 642 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=56160 $D=1
M710 639 631 643 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=60790 $D=1
M711 640 632 644 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=65420 $D=1
M712 641 74 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=51530 $D=1
M713 642 74 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=56160 $D=1
M714 643 74 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=60790 $D=1
M715 644 74 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=65420 $D=1
M716 325 75 641 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=51530 $D=1
M717 326 75 642 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=56160 $D=1
M718 327 75 643 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=60790 $D=1
M719 328 75 644 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=65420 $D=1
M720 645 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=51530 $D=1
M721 646 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=56160 $D=1
M722 647 75 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=60790 $D=1
M723 648 75 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=65420 $D=1
M724 8 76 649 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=51530 $D=1
M725 9 76 650 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=56160 $D=1
M726 10 76 651 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=60790 $D=1
M727 11 76 652 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=65420 $D=1
M728 653 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=51530 $D=1
M729 654 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=56160 $D=1
M730 655 77 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=60790 $D=1
M731 656 77 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=65420 $D=1
M732 657 76 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=51530 $D=1
M733 658 76 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=56160 $D=1
M734 659 76 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=60790 $D=1
M735 660 76 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=65420 $D=1
M736 8 657 1317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=51530 $D=1
M737 9 658 1318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=56160 $D=1
M738 10 659 1319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=60790 $D=1
M739 11 660 1320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=65420 $D=1
M740 661 1317 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=51530 $D=1
M741 662 1318 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=56160 $D=1
M742 663 1319 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=60790 $D=1
M743 664 1320 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=65420 $D=1
M744 657 649 661 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=51530 $D=1
M745 658 650 662 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=56160 $D=1
M746 659 651 663 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=60790 $D=1
M747 660 652 664 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=65420 $D=1
M748 661 77 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=51530 $D=1
M749 662 77 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=56160 $D=1
M750 663 77 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=60790 $D=1
M751 664 77 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=65420 $D=1
M752 325 78 661 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=51530 $D=1
M753 326 78 662 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=56160 $D=1
M754 327 78 663 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=60790 $D=1
M755 328 78 664 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=65420 $D=1
M756 665 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=51530 $D=1
M757 666 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=56160 $D=1
M758 667 78 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=60790 $D=1
M759 668 78 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=65420 $D=1
M760 8 79 669 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=51530 $D=1
M761 9 79 670 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=56160 $D=1
M762 10 79 671 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=60790 $D=1
M763 11 79 672 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=65420 $D=1
M764 673 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=51530 $D=1
M765 674 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=56160 $D=1
M766 675 80 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=60790 $D=1
M767 676 80 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=65420 $D=1
M768 677 79 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=51530 $D=1
M769 678 79 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=56160 $D=1
M770 679 79 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=60790 $D=1
M771 680 79 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=65420 $D=1
M772 8 677 1321 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=51530 $D=1
M773 9 678 1322 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=56160 $D=1
M774 10 679 1323 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=60790 $D=1
M775 11 680 1324 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=65420 $D=1
M776 681 1321 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=51530 $D=1
M777 682 1322 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=56160 $D=1
M778 683 1323 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=60790 $D=1
M779 684 1324 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=65420 $D=1
M780 677 669 681 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=51530 $D=1
M781 678 670 682 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=56160 $D=1
M782 679 671 683 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=60790 $D=1
M783 680 672 684 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=65420 $D=1
M784 681 80 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=51530 $D=1
M785 682 80 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=56160 $D=1
M786 683 80 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=60790 $D=1
M787 684 80 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=65420 $D=1
M788 325 81 681 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=51530 $D=1
M789 326 81 682 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=56160 $D=1
M790 327 81 683 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=60790 $D=1
M791 328 81 684 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=65420 $D=1
M792 685 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=51530 $D=1
M793 686 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=56160 $D=1
M794 687 81 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=60790 $D=1
M795 688 81 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=65420 $D=1
M796 8 82 689 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=51530 $D=1
M797 9 82 690 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=56160 $D=1
M798 10 82 691 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=60790 $D=1
M799 11 82 692 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=65420 $D=1
M800 693 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=51530 $D=1
M801 694 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=56160 $D=1
M802 695 83 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=60790 $D=1
M803 696 83 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=65420 $D=1
M804 697 82 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=51530 $D=1
M805 698 82 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=56160 $D=1
M806 699 82 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=60790 $D=1
M807 700 82 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=65420 $D=1
M808 8 697 1325 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=51530 $D=1
M809 9 698 1326 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=56160 $D=1
M810 10 699 1327 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=60790 $D=1
M811 11 700 1328 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=65420 $D=1
M812 701 1325 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=51530 $D=1
M813 702 1326 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=56160 $D=1
M814 703 1327 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=60790 $D=1
M815 704 1328 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=65420 $D=1
M816 697 689 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=51530 $D=1
M817 698 690 702 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=56160 $D=1
M818 699 691 703 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=60790 $D=1
M819 700 692 704 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=65420 $D=1
M820 701 83 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=51530 $D=1
M821 702 83 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=56160 $D=1
M822 703 83 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=60790 $D=1
M823 704 83 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=65420 $D=1
M824 325 84 701 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=51530 $D=1
M825 326 84 702 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=56160 $D=1
M826 327 84 703 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=60790 $D=1
M827 328 84 704 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=65420 $D=1
M828 705 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=51530 $D=1
M829 706 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=56160 $D=1
M830 707 84 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=60790 $D=1
M831 708 84 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=65420 $D=1
M832 8 85 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=51530 $D=1
M833 9 85 710 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=56160 $D=1
M834 10 85 711 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=60790 $D=1
M835 11 85 712 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=65420 $D=1
M836 713 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=51530 $D=1
M837 714 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=56160 $D=1
M838 715 86 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=60790 $D=1
M839 716 86 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=65420 $D=1
M840 717 85 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=51530 $D=1
M841 718 85 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=56160 $D=1
M842 719 85 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=60790 $D=1
M843 720 85 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=65420 $D=1
M844 8 717 1329 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=51530 $D=1
M845 9 718 1330 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=56160 $D=1
M846 10 719 1331 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=60790 $D=1
M847 11 720 1332 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=65420 $D=1
M848 721 1329 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=51530 $D=1
M849 722 1330 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=56160 $D=1
M850 723 1331 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=60790 $D=1
M851 724 1332 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=65420 $D=1
M852 717 709 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=51530 $D=1
M853 718 710 722 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=56160 $D=1
M854 719 711 723 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=60790 $D=1
M855 720 712 724 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=65420 $D=1
M856 721 86 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=51530 $D=1
M857 722 86 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=56160 $D=1
M858 723 86 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=60790 $D=1
M859 724 86 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=65420 $D=1
M860 325 87 721 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=51530 $D=1
M861 326 87 722 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=56160 $D=1
M862 327 87 723 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=60790 $D=1
M863 328 87 724 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=65420 $D=1
M864 725 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=51530 $D=1
M865 726 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=56160 $D=1
M866 727 87 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=60790 $D=1
M867 728 87 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=65420 $D=1
M868 8 88 729 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=51530 $D=1
M869 9 88 730 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=56160 $D=1
M870 10 88 731 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=60790 $D=1
M871 11 88 732 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=65420 $D=1
M872 733 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=51530 $D=1
M873 734 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=56160 $D=1
M874 735 89 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=60790 $D=1
M875 736 89 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=65420 $D=1
M876 737 88 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=51530 $D=1
M877 738 88 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=56160 $D=1
M878 739 88 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=60790 $D=1
M879 740 88 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=65420 $D=1
M880 8 737 1333 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=51530 $D=1
M881 9 738 1334 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=56160 $D=1
M882 10 739 1335 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=60790 $D=1
M883 11 740 1336 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=65420 $D=1
M884 741 1333 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=51530 $D=1
M885 742 1334 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=56160 $D=1
M886 743 1335 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=60790 $D=1
M887 744 1336 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=65420 $D=1
M888 737 729 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=51530 $D=1
M889 738 730 742 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=56160 $D=1
M890 739 731 743 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=60790 $D=1
M891 740 732 744 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=65420 $D=1
M892 741 89 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=51530 $D=1
M893 742 89 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=56160 $D=1
M894 743 89 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=60790 $D=1
M895 744 89 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=65420 $D=1
M896 325 90 741 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=51530 $D=1
M897 326 90 742 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=56160 $D=1
M898 327 90 743 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=60790 $D=1
M899 328 90 744 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=65420 $D=1
M900 745 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=51530 $D=1
M901 746 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=56160 $D=1
M902 747 90 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=60790 $D=1
M903 748 90 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=65420 $D=1
M904 8 91 749 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=51530 $D=1
M905 9 91 750 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=56160 $D=1
M906 10 91 751 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=60790 $D=1
M907 11 91 752 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=65420 $D=1
M908 753 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=51530 $D=1
M909 754 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=56160 $D=1
M910 755 92 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=60790 $D=1
M911 756 92 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=65420 $D=1
M912 757 91 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=51530 $D=1
M913 758 91 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=56160 $D=1
M914 759 91 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=60790 $D=1
M915 760 91 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=65420 $D=1
M916 8 757 1337 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=51530 $D=1
M917 9 758 1338 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=56160 $D=1
M918 10 759 1339 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=60790 $D=1
M919 11 760 1340 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=65420 $D=1
M920 761 1337 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=51530 $D=1
M921 762 1338 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=56160 $D=1
M922 763 1339 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=60790 $D=1
M923 764 1340 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=65420 $D=1
M924 757 749 761 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=51530 $D=1
M925 758 750 762 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=56160 $D=1
M926 759 751 763 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=60790 $D=1
M927 760 752 764 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=65420 $D=1
M928 761 92 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=51530 $D=1
M929 762 92 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=56160 $D=1
M930 763 92 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=60790 $D=1
M931 764 92 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=65420 $D=1
M932 325 93 761 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=51530 $D=1
M933 326 93 762 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=56160 $D=1
M934 327 93 763 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=60790 $D=1
M935 328 93 764 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=65420 $D=1
M936 765 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=51530 $D=1
M937 766 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=56160 $D=1
M938 767 93 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=60790 $D=1
M939 768 93 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=65420 $D=1
M940 8 94 769 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=51530 $D=1
M941 9 94 770 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=56160 $D=1
M942 10 94 771 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=60790 $D=1
M943 11 94 772 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=65420 $D=1
M944 773 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=51530 $D=1
M945 774 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=56160 $D=1
M946 775 95 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=60790 $D=1
M947 776 95 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=65420 $D=1
M948 777 94 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=51530 $D=1
M949 778 94 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=56160 $D=1
M950 779 94 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=60790 $D=1
M951 780 94 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=65420 $D=1
M952 8 777 1341 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=51530 $D=1
M953 9 778 1342 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=56160 $D=1
M954 10 779 1343 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=60790 $D=1
M955 11 780 1344 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=65420 $D=1
M956 781 1341 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=51530 $D=1
M957 782 1342 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=56160 $D=1
M958 783 1343 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=60790 $D=1
M959 784 1344 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=65420 $D=1
M960 777 769 781 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=51530 $D=1
M961 778 770 782 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=56160 $D=1
M962 779 771 783 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=60790 $D=1
M963 780 772 784 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=65420 $D=1
M964 781 95 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=51530 $D=1
M965 782 95 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=56160 $D=1
M966 783 95 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=60790 $D=1
M967 784 95 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=65420 $D=1
M968 325 96 781 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=51530 $D=1
M969 326 96 782 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=56160 $D=1
M970 327 96 783 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=60790 $D=1
M971 328 96 784 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=65420 $D=1
M972 785 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=51530 $D=1
M973 786 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=56160 $D=1
M974 787 96 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=60790 $D=1
M975 788 96 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=65420 $D=1
M976 8 97 789 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=51530 $D=1
M977 9 97 790 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=56160 $D=1
M978 10 97 791 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=60790 $D=1
M979 11 97 792 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=65420 $D=1
M980 793 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=51530 $D=1
M981 794 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=56160 $D=1
M982 795 98 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=60790 $D=1
M983 796 98 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=65420 $D=1
M984 797 97 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=51530 $D=1
M985 798 97 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=56160 $D=1
M986 799 97 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=60790 $D=1
M987 800 97 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=65420 $D=1
M988 8 797 1345 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=51530 $D=1
M989 9 798 1346 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=56160 $D=1
M990 10 799 1347 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=60790 $D=1
M991 11 800 1348 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=65420 $D=1
M992 801 1345 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=51530 $D=1
M993 802 1346 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=56160 $D=1
M994 803 1347 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=60790 $D=1
M995 804 1348 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=65420 $D=1
M996 797 789 801 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=51530 $D=1
M997 798 790 802 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=56160 $D=1
M998 799 791 803 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=60790 $D=1
M999 800 792 804 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=65420 $D=1
M1000 801 98 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=51530 $D=1
M1001 802 98 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=56160 $D=1
M1002 803 98 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=60790 $D=1
M1003 804 98 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=65420 $D=1
M1004 325 99 801 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=51530 $D=1
M1005 326 99 802 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=56160 $D=1
M1006 327 99 803 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=60790 $D=1
M1007 328 99 804 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=65420 $D=1
M1008 805 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=51530 $D=1
M1009 806 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=56160 $D=1
M1010 807 99 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=60790 $D=1
M1011 808 99 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=65420 $D=1
M1012 8 100 809 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=51530 $D=1
M1013 9 100 810 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=56160 $D=1
M1014 10 100 811 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=60790 $D=1
M1015 11 100 812 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=65420 $D=1
M1016 813 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=51530 $D=1
M1017 814 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=56160 $D=1
M1018 815 101 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=60790 $D=1
M1019 816 101 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=65420 $D=1
M1020 817 100 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=51530 $D=1
M1021 818 100 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=56160 $D=1
M1022 819 100 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=60790 $D=1
M1023 820 100 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=65420 $D=1
M1024 8 817 1349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=51530 $D=1
M1025 9 818 1350 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=56160 $D=1
M1026 10 819 1351 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=60790 $D=1
M1027 11 820 1352 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=65420 $D=1
M1028 821 1349 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=51530 $D=1
M1029 822 1350 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=56160 $D=1
M1030 823 1351 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=60790 $D=1
M1031 824 1352 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=65420 $D=1
M1032 817 809 821 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=51530 $D=1
M1033 818 810 822 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=56160 $D=1
M1034 819 811 823 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=60790 $D=1
M1035 820 812 824 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=65420 $D=1
M1036 821 101 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=51530 $D=1
M1037 822 101 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=56160 $D=1
M1038 823 101 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=60790 $D=1
M1039 824 101 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=65420 $D=1
M1040 325 102 821 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=51530 $D=1
M1041 326 102 822 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=56160 $D=1
M1042 327 102 823 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=60790 $D=1
M1043 328 102 824 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=65420 $D=1
M1044 825 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=51530 $D=1
M1045 826 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=56160 $D=1
M1046 827 102 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=60790 $D=1
M1047 828 102 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=65420 $D=1
M1048 8 103 829 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=51530 $D=1
M1049 9 103 830 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=56160 $D=1
M1050 10 103 831 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=60790 $D=1
M1051 11 103 832 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=65420 $D=1
M1052 833 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=51530 $D=1
M1053 834 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=56160 $D=1
M1054 835 104 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=60790 $D=1
M1055 836 104 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=65420 $D=1
M1056 837 103 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=51530 $D=1
M1057 838 103 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=56160 $D=1
M1058 839 103 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=60790 $D=1
M1059 840 103 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=65420 $D=1
M1060 8 837 1353 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=51530 $D=1
M1061 9 838 1354 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=56160 $D=1
M1062 10 839 1355 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=60790 $D=1
M1063 11 840 1356 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=65420 $D=1
M1064 841 1353 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=51530 $D=1
M1065 842 1354 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=56160 $D=1
M1066 843 1355 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=60790 $D=1
M1067 844 1356 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=65420 $D=1
M1068 837 829 841 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=51530 $D=1
M1069 838 830 842 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=56160 $D=1
M1070 839 831 843 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=60790 $D=1
M1071 840 832 844 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=65420 $D=1
M1072 841 104 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=51530 $D=1
M1073 842 104 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=56160 $D=1
M1074 843 104 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=60790 $D=1
M1075 844 104 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=65420 $D=1
M1076 325 105 841 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=51530 $D=1
M1077 326 105 842 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=56160 $D=1
M1078 327 105 843 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=60790 $D=1
M1079 328 105 844 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=65420 $D=1
M1080 845 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=51530 $D=1
M1081 846 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=56160 $D=1
M1082 847 105 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=60790 $D=1
M1083 848 105 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=65420 $D=1
M1084 8 106 849 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=51530 $D=1
M1085 9 106 850 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=56160 $D=1
M1086 10 106 851 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=60790 $D=1
M1087 11 106 852 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=65420 $D=1
M1088 853 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=51530 $D=1
M1089 854 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=56160 $D=1
M1090 855 107 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=60790 $D=1
M1091 856 107 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=65420 $D=1
M1092 857 106 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=51530 $D=1
M1093 858 106 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=56160 $D=1
M1094 859 106 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=60790 $D=1
M1095 860 106 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=65420 $D=1
M1096 8 857 1357 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=51530 $D=1
M1097 9 858 1358 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=56160 $D=1
M1098 10 859 1359 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=60790 $D=1
M1099 11 860 1360 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=65420 $D=1
M1100 861 1357 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=51530 $D=1
M1101 862 1358 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=56160 $D=1
M1102 863 1359 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=60790 $D=1
M1103 864 1360 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=65420 $D=1
M1104 857 849 861 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=51530 $D=1
M1105 858 850 862 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=56160 $D=1
M1106 859 851 863 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=60790 $D=1
M1107 860 852 864 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=65420 $D=1
M1108 861 107 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=51530 $D=1
M1109 862 107 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=56160 $D=1
M1110 863 107 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=60790 $D=1
M1111 864 107 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=65420 $D=1
M1112 325 108 861 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=51530 $D=1
M1113 326 108 862 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=56160 $D=1
M1114 327 108 863 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=60790 $D=1
M1115 328 108 864 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=65420 $D=1
M1116 865 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=51530 $D=1
M1117 866 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=56160 $D=1
M1118 867 108 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=60790 $D=1
M1119 868 108 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=65420 $D=1
M1120 8 109 869 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=51530 $D=1
M1121 9 109 870 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=56160 $D=1
M1122 10 109 871 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=60790 $D=1
M1123 11 109 872 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=65420 $D=1
M1124 873 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=51530 $D=1
M1125 874 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=56160 $D=1
M1126 875 110 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=60790 $D=1
M1127 876 110 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=65420 $D=1
M1128 877 109 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=51530 $D=1
M1129 878 109 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=56160 $D=1
M1130 879 109 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=60790 $D=1
M1131 880 109 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=65420 $D=1
M1132 8 877 1361 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=51530 $D=1
M1133 9 878 1362 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=56160 $D=1
M1134 10 879 1363 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=60790 $D=1
M1135 11 880 1364 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=65420 $D=1
M1136 881 1361 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=51530 $D=1
M1137 882 1362 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=56160 $D=1
M1138 883 1363 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=60790 $D=1
M1139 884 1364 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=65420 $D=1
M1140 877 869 881 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=51530 $D=1
M1141 878 870 882 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=56160 $D=1
M1142 879 871 883 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=60790 $D=1
M1143 880 872 884 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=65420 $D=1
M1144 881 110 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=51530 $D=1
M1145 882 110 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=56160 $D=1
M1146 883 110 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=60790 $D=1
M1147 884 110 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=65420 $D=1
M1148 325 111 881 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=51530 $D=1
M1149 326 111 882 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=56160 $D=1
M1150 327 111 883 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=60790 $D=1
M1151 328 111 884 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=65420 $D=1
M1152 885 111 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=51530 $D=1
M1153 886 111 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=56160 $D=1
M1154 887 111 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=60790 $D=1
M1155 888 111 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=65420 $D=1
M1156 8 112 889 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=51530 $D=1
M1157 9 112 890 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=56160 $D=1
M1158 10 112 891 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=60790 $D=1
M1159 11 112 892 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=65420 $D=1
M1160 893 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=51530 $D=1
M1161 894 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=56160 $D=1
M1162 895 113 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=60790 $D=1
M1163 896 113 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=65420 $D=1
M1164 897 112 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=51530 $D=1
M1165 898 112 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=56160 $D=1
M1166 899 112 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=60790 $D=1
M1167 900 112 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=65420 $D=1
M1168 8 897 1365 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=51530 $D=1
M1169 9 898 1366 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=56160 $D=1
M1170 10 899 1367 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=60790 $D=1
M1171 11 900 1368 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=65420 $D=1
M1172 901 1365 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=51530 $D=1
M1173 902 1366 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=56160 $D=1
M1174 903 1367 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=60790 $D=1
M1175 904 1368 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=65420 $D=1
M1176 897 889 901 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=51530 $D=1
M1177 898 890 902 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=56160 $D=1
M1178 899 891 903 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=60790 $D=1
M1179 900 892 904 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=65420 $D=1
M1180 901 113 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=51530 $D=1
M1181 902 113 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=56160 $D=1
M1182 903 113 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=60790 $D=1
M1183 904 113 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=65420 $D=1
M1184 325 116 901 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=51530 $D=1
M1185 326 116 902 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=56160 $D=1
M1186 327 116 903 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=60790 $D=1
M1187 328 116 904 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=65420 $D=1
M1188 905 116 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=51530 $D=1
M1189 906 116 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=56160 $D=1
M1190 907 116 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=60790 $D=1
M1191 908 116 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=65420 $D=1
M1192 8 117 909 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=51530 $D=1
M1193 9 117 910 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=56160 $D=1
M1194 10 117 911 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=60790 $D=1
M1195 11 117 912 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=65420 $D=1
M1196 913 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=51530 $D=1
M1197 914 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=56160 $D=1
M1198 915 118 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=60790 $D=1
M1199 916 118 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=65420 $D=1
M1200 917 117 297 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=51530 $D=1
M1201 918 117 298 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=56160 $D=1
M1202 919 117 299 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=60790 $D=1
M1203 920 117 300 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=65420 $D=1
M1204 8 917 1369 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=51530 $D=1
M1205 9 918 1370 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=56160 $D=1
M1206 10 919 1371 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=60790 $D=1
M1207 11 920 1372 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=65420 $D=1
M1208 921 1369 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=51530 $D=1
M1209 922 1370 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=56160 $D=1
M1210 923 1371 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=60790 $D=1
M1211 924 1372 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=65420 $D=1
M1212 917 909 921 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=51530 $D=1
M1213 918 910 922 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=56160 $D=1
M1214 919 911 923 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=60790 $D=1
M1215 920 912 924 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=65420 $D=1
M1216 921 118 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=51530 $D=1
M1217 922 118 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=56160 $D=1
M1218 923 118 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=60790 $D=1
M1219 924 118 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=65420 $D=1
M1220 325 122 921 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=51530 $D=1
M1221 326 122 922 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=56160 $D=1
M1222 327 122 923 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=60790 $D=1
M1223 328 122 924 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=65420 $D=1
M1224 925 122 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=51530 $D=1
M1225 926 122 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=56160 $D=1
M1226 927 122 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=60790 $D=1
M1227 928 122 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=65420 $D=1
M1228 8 123 929 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=51530 $D=1
M1229 9 123 930 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=56160 $D=1
M1230 10 123 931 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=60790 $D=1
M1231 11 123 932 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=65420 $D=1
M1232 933 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=51530 $D=1
M1233 934 124 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=56160 $D=1
M1234 935 124 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=60790 $D=1
M1235 936 124 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=65420 $D=1
M1236 8 124 317 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=51530 $D=1
M1237 9 124 318 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=56160 $D=1
M1238 10 124 319 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=60790 $D=1
M1239 11 124 320 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=65420 $D=1
M1240 325 123 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=51530 $D=1
M1241 326 123 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=56160 $D=1
M1242 327 123 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=60790 $D=1
M1243 328 123 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=65420 $D=1
M1244 8 941 937 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=51530 $D=1
M1245 9 942 938 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=56160 $D=1
M1246 10 943 939 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=60790 $D=1
M1247 11 944 940 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=65420 $D=1
M1248 941 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=51530 $D=1
M1249 942 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=56160 $D=1
M1250 943 126 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=60790 $D=1
M1251 944 126 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=65420 $D=1
M1252 1373 317 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=51530 $D=1
M1253 1374 318 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=56160 $D=1
M1254 1375 319 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=60790 $D=1
M1255 1376 320 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=65420 $D=1
M1256 945 937 1373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=51530 $D=1
M1257 946 938 1374 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=56160 $D=1
M1258 947 939 1375 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=60790 $D=1
M1259 948 940 1376 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=65420 $D=1
M1260 8 945 949 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=51530 $D=1
M1261 9 946 950 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=56160 $D=1
M1262 10 947 951 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=60790 $D=1
M1263 11 948 952 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=65420 $D=1
M1264 1377 949 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=51530 $D=1
M1265 1378 950 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=56160 $D=1
M1266 1379 951 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=60790 $D=1
M1267 1380 952 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=65420 $D=1
M1268 945 941 1377 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=51530 $D=1
M1269 946 942 1378 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=56160 $D=1
M1270 947 943 1379 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=60790 $D=1
M1271 948 944 1380 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=65420 $D=1
M1272 8 957 953 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=51530 $D=1
M1273 9 958 954 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=56160 $D=1
M1274 10 959 955 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=60790 $D=1
M1275 11 960 956 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=65420 $D=1
M1276 957 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=51530 $D=1
M1277 958 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=56160 $D=1
M1278 959 126 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=60790 $D=1
M1279 960 126 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=65420 $D=1
M1280 1381 325 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=51530 $D=1
M1281 1382 326 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=56160 $D=1
M1282 1383 327 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=60790 $D=1
M1283 1384 328 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=65420 $D=1
M1284 961 953 1381 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=51530 $D=1
M1285 962 954 1382 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=56160 $D=1
M1286 963 955 1383 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=60790 $D=1
M1287 964 956 1384 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=65420 $D=1
M1288 8 961 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=51530 $D=1
M1289 9 962 128 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=56160 $D=1
M1290 10 963 129 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=60790 $D=1
M1291 11 964 130 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=65420 $D=1
M1292 1385 127 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=51530 $D=1
M1293 1386 128 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=56160 $D=1
M1294 1387 129 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=60790 $D=1
M1295 1388 130 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=65420 $D=1
M1296 961 957 1385 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=51530 $D=1
M1297 962 958 1386 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=56160 $D=1
M1298 963 959 1387 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=60790 $D=1
M1299 964 960 1388 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=65420 $D=1
M1300 965 131 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=51530 $D=1
M1301 966 131 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=56160 $D=1
M1302 967 131 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=60790 $D=1
M1303 968 131 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=65420 $D=1
M1304 969 965 949 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=51530 $D=1
M1305 970 966 950 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=56160 $D=1
M1306 971 967 951 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=60790 $D=1
M1307 972 968 952 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=65420 $D=1
M1308 132 131 969 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=51530 $D=1
M1309 132 131 970 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=56160 $D=1
M1310 132 131 971 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=60790 $D=1
M1311 132 131 972 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=65420 $D=1
M1312 973 133 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=51530 $D=1
M1313 974 133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=56160 $D=1
M1314 975 133 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=60790 $D=1
M1315 976 133 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=65420 $D=1
M1316 977 973 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=51530 $D=1
M1317 978 974 128 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=56160 $D=1
M1318 979 975 129 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=60790 $D=1
M1319 980 976 130 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=65420 $D=1
M1320 1389 133 977 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=51530 $D=1
M1321 1390 133 978 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=56160 $D=1
M1322 1391 133 979 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=60790 $D=1
M1323 1392 133 980 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=65420 $D=1
M1324 8 127 1389 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=51530 $D=1
M1325 9 128 1390 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=56160 $D=1
M1326 10 129 1391 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=60790 $D=1
M1327 11 130 1392 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=65420 $D=1
M1328 981 134 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=51530 $D=1
M1329 982 134 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=56160 $D=1
M1330 983 134 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=60790 $D=1
M1331 984 134 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=65420 $D=1
M1332 985 981 977 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=51530 $D=1
M1333 986 982 978 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=56160 $D=1
M1334 987 983 979 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=60790 $D=1
M1335 988 984 980 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=65420 $D=1
M1336 15 134 985 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=51530 $D=1
M1337 16 134 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=56160 $D=1
M1338 17 134 987 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=60790 $D=1
M1339 18 134 988 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=65420 $D=1
M1340 992 989 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=51530 $D=1
M1341 993 990 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=56160 $D=1
M1342 994 991 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=60790 $D=1
M1343 995 135 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=65420 $D=1
M1344 8 1000 996 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=51530 $D=1
M1345 9 1001 997 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=56160 $D=1
M1346 10 1002 998 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=60790 $D=1
M1347 11 1003 999 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=65420 $D=1
M1348 1004 969 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=51530 $D=1
M1349 1005 970 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=56160 $D=1
M1350 1006 971 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=60790 $D=1
M1351 1007 972 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=65420 $D=1
M1352 1000 1004 989 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=51530 $D=1
M1353 1001 1005 990 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=56160 $D=1
M1354 1002 1006 991 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=60790 $D=1
M1355 1003 1007 135 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=65420 $D=1
M1356 992 969 1000 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=51530 $D=1
M1357 993 970 1001 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=56160 $D=1
M1358 994 971 1002 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=60790 $D=1
M1359 995 972 1003 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=65420 $D=1
M1360 1008 996 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=51530 $D=1
M1361 1009 997 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=56160 $D=1
M1362 1010 998 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=60790 $D=1
M1363 1011 999 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=65420 $D=1
M1364 136 1008 985 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=51530 $D=1
M1365 989 1009 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=56160 $D=1
M1366 990 1010 987 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=60790 $D=1
M1367 991 1011 988 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=65420 $D=1
M1368 969 996 136 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=51530 $D=1
M1369 970 997 989 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=56160 $D=1
M1370 971 998 990 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=60790 $D=1
M1371 972 999 991 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=65420 $D=1
M1372 1012 136 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=51530 $D=1
M1373 1013 989 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=56160 $D=1
M1374 1014 990 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=60790 $D=1
M1375 1015 991 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=65420 $D=1
M1376 1016 996 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=51530 $D=1
M1377 1017 997 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=56160 $D=1
M1378 1018 998 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=60790 $D=1
M1379 1019 999 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=65420 $D=1
M1380 1020 1016 1012 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=51530 $D=1
M1381 1021 1017 1013 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=56160 $D=1
M1382 1022 1018 1014 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=60790 $D=1
M1383 1023 1019 1015 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=65420 $D=1
M1384 985 996 1020 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=51530 $D=1
M1385 986 997 1021 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=56160 $D=1
M1386 987 998 1022 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=60790 $D=1
M1387 988 999 1023 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=65420 $D=1
M1388 1024 969 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=51530 $D=1
M1389 1025 970 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=56160 $D=1
M1390 1026 971 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=60790 $D=1
M1391 1027 972 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=65420 $D=1
M1392 8 985 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=51530 $D=1
M1393 9 986 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=56160 $D=1
M1394 10 987 1026 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=60790 $D=1
M1395 11 988 1027 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=65420 $D=1
M1396 1028 1020 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=51530 $D=1
M1397 1029 1021 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=56160 $D=1
M1398 1030 1022 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=60790 $D=1
M1399 1031 1023 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=65420 $D=1
M1400 1429 969 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=51530 $D=1
M1401 1430 970 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=56160 $D=1
M1402 1431 971 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=60790 $D=1
M1403 1432 972 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=65420 $D=1
M1404 1032 985 1429 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=51530 $D=1
M1405 1033 986 1430 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=56160 $D=1
M1406 1034 987 1431 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=60790 $D=1
M1407 1035 988 1432 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=65420 $D=1
M1408 1433 969 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=51530 $D=1
M1409 1434 970 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=56160 $D=1
M1410 1435 971 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=60790 $D=1
M1411 1436 972 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=65420 $D=1
M1412 1036 985 1433 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=51530 $D=1
M1413 1037 986 1434 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=56160 $D=1
M1414 1038 987 1435 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=60790 $D=1
M1415 1039 988 1436 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=65420 $D=1
M1416 1044 969 1040 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=51530 $D=1
M1417 1045 970 1041 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=56160 $D=1
M1418 1046 971 1042 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=60790 $D=1
M1419 1047 972 1043 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=65420 $D=1
M1420 1040 985 1044 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=51530 $D=1
M1421 1041 986 1045 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=56160 $D=1
M1422 1042 987 1046 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=60790 $D=1
M1423 1043 988 1047 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=65420 $D=1
M1424 8 1036 1040 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=51530 $D=1
M1425 9 1037 1041 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=56160 $D=1
M1426 10 1038 1042 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=60790 $D=1
M1427 11 1039 1043 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=65420 $D=1
M1428 1048 140 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=51530 $D=1
M1429 1049 140 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=56160 $D=1
M1430 1050 140 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=60790 $D=1
M1431 1051 140 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=65420 $D=1
M1432 1052 1048 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=51530 $D=1
M1433 1053 1049 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=56160 $D=1
M1434 1054 1050 1026 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=60790 $D=1
M1435 1055 1051 1027 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=65420 $D=1
M1436 1032 140 1052 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=51530 $D=1
M1437 1033 140 1053 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=56160 $D=1
M1438 1034 140 1054 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=60790 $D=1
M1439 1035 140 1055 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=65420 $D=1
M1440 1056 1048 1028 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=51530 $D=1
M1441 1057 1049 1029 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=56160 $D=1
M1442 1058 1050 1030 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=60790 $D=1
M1443 1059 1051 1031 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=65420 $D=1
M1444 1044 140 1056 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=51530 $D=1
M1445 1045 140 1057 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=56160 $D=1
M1446 1046 140 1058 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=60790 $D=1
M1447 1047 140 1059 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=65420 $D=1
M1448 1060 141 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=51530 $D=1
M1449 1061 141 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=56160 $D=1
M1450 1062 141 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=60790 $D=1
M1451 1063 141 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=65420 $D=1
M1452 1064 1060 1056 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=51530 $D=1
M1453 1065 1061 1057 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=56160 $D=1
M1454 1066 1062 1058 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=60790 $D=1
M1455 1067 1063 1059 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=65420 $D=1
M1456 1052 141 1064 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=51530 $D=1
M1457 1053 141 1065 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=56160 $D=1
M1458 1054 141 1066 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=60790 $D=1
M1459 1055 141 1067 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=65420 $D=1
M1460 19 1064 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=51530 $D=1
M1461 20 1065 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=56160 $D=1
M1462 21 1066 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=60790 $D=1
M1463 22 1067 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=65420 $D=1
M1464 1068 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=51530 $D=1
M1465 1069 142 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=56160 $D=1
M1466 1070 142 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=60790 $D=1
M1467 1071 142 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=65420 $D=1
M1468 1072 1068 143 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=51530 $D=1
M1469 1073 1069 144 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=56160 $D=1
M1470 1074 1070 145 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=60790 $D=1
M1471 1075 1071 146 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=65420 $D=1
M1472 147 142 1072 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=51530 $D=1
M1473 148 142 1073 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=56160 $D=1
M1474 143 142 1074 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=60790 $D=1
M1475 144 142 1075 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=65420 $D=1
M1476 1076 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=51530 $D=1
M1477 1077 142 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=56160 $D=1
M1478 1078 142 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=60790 $D=1
M1479 1079 142 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=65420 $D=1
M1480 1080 1076 149 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=51530 $D=1
M1481 1081 1077 150 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=56160 $D=1
M1482 1082 1078 151 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=60790 $D=1
M1483 1083 1079 152 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=65420 $D=1
M1484 153 142 1080 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=51530 $D=1
M1485 154 142 1081 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=56160 $D=1
M1486 155 142 1082 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=60790 $D=1
M1487 156 142 1083 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=65420 $D=1
M1488 1084 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=51530 $D=1
M1489 1085 142 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=56160 $D=1
M1490 1086 142 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=60790 $D=1
M1491 1087 142 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=65420 $D=1
M1492 1088 1084 137 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=51530 $D=1
M1493 1089 1085 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=56160 $D=1
M1494 1090 1086 138 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=60790 $D=1
M1495 1091 1087 157 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=65420 $D=1
M1496 158 142 1088 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=51530 $D=1
M1497 120 142 1089 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=56160 $D=1
M1498 121 142 1090 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=60790 $D=1
M1499 125 142 1091 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=65420 $D=1
M1500 1092 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=51530 $D=1
M1501 1093 142 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=56160 $D=1
M1502 1094 142 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=60790 $D=1
M1503 1095 142 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=65420 $D=1
M1504 1096 1092 159 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=51530 $D=1
M1505 1097 1093 160 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=56160 $D=1
M1506 1098 1094 161 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=60790 $D=1
M1507 1099 1095 162 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=65420 $D=1
M1508 163 142 1096 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=51530 $D=1
M1509 164 142 1097 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=56160 $D=1
M1510 165 142 1098 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=60790 $D=1
M1511 166 142 1099 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=65420 $D=1
M1512 1100 142 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=51530 $D=1
M1513 1101 142 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=56160 $D=1
M1514 1102 142 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=60790 $D=1
M1515 1103 142 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=65420 $D=1
M1516 1104 1100 167 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=51530 $D=1
M1517 1105 1101 168 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=56160 $D=1
M1518 1106 1102 169 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=60790 $D=1
M1519 1107 1103 170 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=65420 $D=1
M1520 171 142 1104 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=51530 $D=1
M1521 171 142 1105 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=56160 $D=1
M1522 171 142 1106 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=60790 $D=1
M1523 171 142 1107 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=65420 $D=1
M1524 8 969 1393 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=51530 $D=1
M1525 9 970 1394 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=56160 $D=1
M1526 10 971 1395 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=60790 $D=1
M1527 11 972 1396 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=65420 $D=1
M1528 148 1393 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=51530 $D=1
M1529 143 1394 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=56160 $D=1
M1530 144 1395 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=60790 $D=1
M1531 145 1396 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=65420 $D=1
M1532 1108 172 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=51530 $D=1
M1533 1109 172 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=56160 $D=1
M1534 1110 172 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=60790 $D=1
M1535 1111 172 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=65420 $D=1
M1536 155 1108 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=51530 $D=1
M1537 156 1109 143 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=56160 $D=1
M1538 149 1110 144 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=60790 $D=1
M1539 150 1111 145 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=65420 $D=1
M1540 1072 172 155 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=51530 $D=1
M1541 1073 172 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=56160 $D=1
M1542 1074 172 149 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=60790 $D=1
M1543 1075 172 150 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=65420 $D=1
M1544 1112 173 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=51530 $D=1
M1545 1113 173 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=56160 $D=1
M1546 1114 173 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=60790 $D=1
M1547 1115 173 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=65420 $D=1
M1548 174 1112 155 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=51530 $D=1
M1549 114 1113 156 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=56160 $D=1
M1550 115 1114 149 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=60790 $D=1
M1551 119 1115 150 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=65420 $D=1
M1552 1080 173 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=51530 $D=1
M1553 1081 173 114 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=56160 $D=1
M1554 1082 173 115 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=60790 $D=1
M1555 1083 173 119 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=65420 $D=1
M1556 1116 175 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=51530 $D=1
M1557 1117 175 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=56160 $D=1
M1558 1118 175 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=60790 $D=1
M1559 1119 175 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=65420 $D=1
M1560 174 1116 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=51530 $D=1
M1561 114 1117 114 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=56160 $D=1
M1562 115 1118 115 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=60790 $D=1
M1563 119 1119 119 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=65420 $D=1
M1564 1088 175 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=51530 $D=1
M1565 1089 175 114 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=56160 $D=1
M1566 1090 175 115 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=60790 $D=1
M1567 1091 175 119 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=65420 $D=1
M1568 1120 176 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=51530 $D=1
M1569 1121 176 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=56160 $D=1
M1570 1122 176 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=60790 $D=1
M1571 1123 176 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=65420 $D=1
M1572 177 1120 174 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=51530 $D=1
M1573 178 1121 114 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=56160 $D=1
M1574 179 1122 115 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=60790 $D=1
M1575 180 1123 119 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=65420 $D=1
M1576 1096 176 177 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=51530 $D=1
M1577 1097 176 178 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=56160 $D=1
M1578 1098 176 179 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=60790 $D=1
M1579 1099 176 180 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=65420 $D=1
M1580 1124 181 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=51530 $D=1
M1581 1125 181 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=56160 $D=1
M1582 1126 181 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=60790 $D=1
M1583 1127 181 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=65420 $D=1
M1584 269 1124 177 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=51530 $D=1
M1585 270 1125 178 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=56160 $D=1
M1586 271 1126 179 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=60790 $D=1
M1587 272 1127 180 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=65420 $D=1
M1588 1104 181 269 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=51530 $D=1
M1589 1105 181 270 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=56160 $D=1
M1590 1106 181 271 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=60790 $D=1
M1591 1107 181 272 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=65420 $D=1
M1592 1128 182 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=51530 $D=1
M1593 1129 182 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=56160 $D=1
M1594 1130 182 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=60790 $D=1
M1595 1131 182 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=65420 $D=1
M1596 1132 1128 127 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=51530 $D=1
M1597 1133 1129 128 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=56160 $D=1
M1598 1134 1130 129 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=60790 $D=1
M1599 1135 1131 130 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=65420 $D=1
M1600 15 182 1132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=51530 $D=1
M1601 16 182 1133 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=56160 $D=1
M1602 17 182 1134 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=60790 $D=1
M1603 18 182 1135 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=65420 $D=1
M1604 1437 949 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=51530 $D=1
M1605 1438 950 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=56160 $D=1
M1606 1439 951 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=60790 $D=1
M1607 1440 952 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=65420 $D=1
M1608 1136 1132 1437 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=51530 $D=1
M1609 1137 1133 1438 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=56160 $D=1
M1610 1138 1134 1439 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=60790 $D=1
M1611 1139 1135 1440 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=65420 $D=1
M1612 1144 949 1140 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=51530 $D=1
M1613 1145 950 1141 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=56160 $D=1
M1614 1146 951 1142 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=60790 $D=1
M1615 1147 952 1143 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=65420 $D=1
M1616 1140 1132 1144 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=51530 $D=1
M1617 1141 1133 1145 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=56160 $D=1
M1618 1142 1134 1146 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=60790 $D=1
M1619 1143 1135 1147 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=65420 $D=1
M1620 8 1136 1140 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=51530 $D=1
M1621 9 1137 1141 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=56160 $D=1
M1622 10 1138 1142 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=60790 $D=1
M1623 11 1139 1143 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=65420 $D=1
M1624 1441 183 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=51530 $D=1
M1625 1442 1148 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=56160 $D=1
M1626 1443 1149 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=60790 $D=1
M1627 1444 1150 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=65420 $D=1
M1628 1397 1144 1441 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=51530 $D=1
M1629 1398 1145 1442 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=56160 $D=1
M1630 1399 1146 1443 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=60790 $D=1
M1631 1400 1147 1444 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=65420 $D=1
M1632 1148 1397 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=51530 $D=1
M1633 1149 1398 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=56160 $D=1
M1634 1150 1399 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=60790 $D=1
M1635 184 1400 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=65420 $D=1
M1636 1151 949 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=51530 $D=1
M1637 1152 950 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=56160 $D=1
M1638 1153 951 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=60790 $D=1
M1639 1154 952 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=65420 $D=1
M1640 8 1155 1151 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=51530 $D=1
M1641 9 1156 1152 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=56160 $D=1
M1642 10 1157 1153 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=60790 $D=1
M1643 11 1158 1154 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=65420 $D=1
M1644 1155 1132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=51530 $D=1
M1645 1156 1133 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=56160 $D=1
M1646 1157 1134 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=60790 $D=1
M1647 1158 1135 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=65420 $D=1
M1648 1445 1151 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=51530 $D=1
M1649 1446 1152 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=56160 $D=1
M1650 1447 1153 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=60790 $D=1
M1651 1448 1154 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=65420 $D=1
M1652 1159 183 1445 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=51530 $D=1
M1653 1160 1148 1446 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=56160 $D=1
M1654 1161 1149 1447 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=60790 $D=1
M1655 1162 1150 1448 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=65420 $D=1
M1656 1166 185 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=51530 $D=1
M1657 1167 1163 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=56160 $D=1
M1658 1168 1164 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=60790 $D=1
M1659 1169 1165 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=65420 $D=1
M1660 1449 1159 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=51530 $D=1
M1661 1450 1160 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=56160 $D=1
M1662 1451 1161 10 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=60790 $D=1
M1663 1452 1162 11 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=65420 $D=1
M1664 1163 1166 1449 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=51530 $D=1
M1665 1164 1167 1450 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=56160 $D=1
M1666 1165 1168 1451 10 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=60790 $D=1
M1667 186 1169 1452 11 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=65420 $D=1
M1668 1173 1170 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=51530 $D=1
M1669 1174 1171 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=56160 $D=1
M1670 1175 1172 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=60790 $D=1
M1671 1176 187 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=65420 $D=1
M1672 8 1181 1177 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=51530 $D=1
M1673 9 1182 1178 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=56160 $D=1
M1674 10 1183 1179 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=60790 $D=1
M1675 11 1184 1180 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=65420 $D=1
M1676 1185 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=51530 $D=1
M1677 1186 132 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=56160 $D=1
M1678 1187 132 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=60790 $D=1
M1679 1188 132 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=65420 $D=1
M1680 1181 1185 1170 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=51530 $D=1
M1681 1182 1186 1171 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=56160 $D=1
M1682 1183 1187 1172 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=60790 $D=1
M1683 1184 1188 187 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=65420 $D=1
M1684 1173 132 1181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=51530 $D=1
M1685 1174 132 1182 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=56160 $D=1
M1686 1175 132 1183 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=60790 $D=1
M1687 1176 132 1184 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=65420 $D=1
M1688 1189 1177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=51530 $D=1
M1689 1190 1178 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=56160 $D=1
M1690 1191 1179 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=60790 $D=1
M1691 1192 1180 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=65420 $D=1
M1692 188 1189 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=51530 $D=1
M1693 1170 1190 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=56160 $D=1
M1694 1171 1191 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=60790 $D=1
M1695 1172 1192 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=65420 $D=1
M1696 132 1177 188 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=51530 $D=1
M1697 132 1178 1170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=56160 $D=1
M1698 132 1179 1171 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=60790 $D=1
M1699 132 1180 1172 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=65420 $D=1
M1700 1193 188 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=51530 $D=1
M1701 1194 1170 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=56160 $D=1
M1702 1195 1171 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=60790 $D=1
M1703 1196 1172 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=65420 $D=1
M1704 1197 1177 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=51530 $D=1
M1705 1198 1178 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=56160 $D=1
M1706 1199 1179 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=60790 $D=1
M1707 1200 1180 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=65420 $D=1
M1708 273 1197 1193 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=51530 $D=1
M1709 274 1198 1194 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=56160 $D=1
M1710 275 1199 1195 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=60790 $D=1
M1711 276 1200 1196 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=65420 $D=1
M1712 8 1177 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=51530 $D=1
M1713 9 1178 274 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=56160 $D=1
M1714 10 1179 275 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=60790 $D=1
M1715 11 1180 276 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=65420 $D=1
M1716 1201 189 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=51530 $D=1
M1717 1202 189 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=56160 $D=1
M1718 1203 189 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=60790 $D=1
M1719 1204 189 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=65420 $D=1
M1720 1205 1201 273 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=51530 $D=1
M1721 1206 1202 274 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=56160 $D=1
M1722 1207 1203 275 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=60790 $D=1
M1723 1208 1204 276 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=65420 $D=1
M1724 19 189 1205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=51530 $D=1
M1725 20 189 1206 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=56160 $D=1
M1726 21 189 1207 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=60790 $D=1
M1727 22 189 1208 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=65420 $D=1
M1728 1209 190 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=51530 $D=1
M1729 1210 190 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=56160 $D=1
M1730 1211 190 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=60790 $D=1
M1731 1212 190 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=65420 $D=1
M1732 190 1209 1205 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=51530 $D=1
M1733 190 1210 1206 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=56160 $D=1
M1734 190 1211 1207 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=60790 $D=1
M1735 190 1212 1208 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=65420 $D=1
M1736 8 190 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=51530 $D=1
M1737 9 190 190 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=56160 $D=1
M1738 10 190 190 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=60790 $D=1
M1739 11 190 190 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=65420 $D=1
M1740 1213 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=51530 $D=1
M1741 1214 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=56160 $D=1
M1742 1215 126 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=60790 $D=1
M1743 1216 126 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=65420 $D=1
M1744 8 1213 1217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=51530 $D=1
M1745 9 1214 1218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=56160 $D=1
M1746 10 1215 1219 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=60790 $D=1
M1747 11 1216 1220 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=65420 $D=1
M1748 1221 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=51530 $D=1
M1749 1222 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=56160 $D=1
M1750 1223 126 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=60790 $D=1
M1751 1224 126 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=65420 $D=1
M1752 1225 1213 190 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=51530 $D=1
M1753 1226 1214 190 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=56160 $D=1
M1754 1227 1215 190 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=60790 $D=1
M1755 1228 1216 190 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=65420 $D=1
M1756 8 1225 1401 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=51530 $D=1
M1757 9 1226 1402 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=56160 $D=1
M1758 10 1227 1403 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=60790 $D=1
M1759 11 1228 1404 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=65420 $D=1
M1760 1229 1401 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=51530 $D=1
M1761 1230 1402 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=56160 $D=1
M1762 1231 1403 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=60790 $D=1
M1763 1232 1404 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=65420 $D=1
M1764 1225 1217 1229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=51530 $D=1
M1765 1226 1218 1230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=56160 $D=1
M1766 1227 1219 1231 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=60790 $D=1
M1767 1228 1220 1232 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=65420 $D=1
M1768 1233 126 1229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=51530 $D=1
M1769 1234 126 1230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=56160 $D=1
M1770 1235 126 1231 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=60790 $D=1
M1771 1236 126 1232 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=65420 $D=1
M1772 8 1241 1237 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=51530 $D=1
M1773 9 1242 1238 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=56160 $D=1
M1774 10 1243 1239 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=60790 $D=1
M1775 11 1244 1240 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=65420 $D=1
M1776 1241 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=51530 $D=1
M1777 1242 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=56160 $D=1
M1778 1243 126 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=60790 $D=1
M1779 1244 126 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=65420 $D=1
M1780 1405 1233 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=51530 $D=1
M1781 1406 1234 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=56160 $D=1
M1782 1407 1235 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=60790 $D=1
M1783 1408 1236 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=65420 $D=1
M1784 1245 1237 1405 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=51530 $D=1
M1785 1246 1238 1406 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=56160 $D=1
M1786 1247 1239 1407 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=60790 $D=1
M1787 1248 1240 1408 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=65420 $D=1
M1788 8 1245 132 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=51530 $D=1
M1789 9 1246 132 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=56160 $D=1
M1790 10 1247 132 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=60790 $D=1
M1791 11 1248 132 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=65420 $D=1
M1792 1409 132 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=51530 $D=1
M1793 1410 132 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=56160 $D=1
M1794 1411 132 10 10 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=60790 $D=1
M1795 1412 132 11 11 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=65420 $D=1
M1796 1245 1241 1409 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=51530 $D=1
M1797 1246 1242 1410 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=56160 $D=1
M1798 1247 1243 1411 10 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=60790 $D=1
M1799 1248 1244 1412 11 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=65420 $D=1
M1800 221 1 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=52780 $D=0
M1801 222 1 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=57410 $D=0
M1802 223 1 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=62040 $D=0
M1803 224 1 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=66670 $D=0
M1804 225 1 2 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=52780 $D=0
M1805 226 1 3 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=57410 $D=0
M1806 227 1 4 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=62040 $D=0
M1807 228 1 5 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=66670 $D=0
M1808 8 221 225 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=52780 $D=0
M1809 9 222 226 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=57410 $D=0
M1810 10 223 227 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=62040 $D=0
M1811 11 224 228 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=66670 $D=0
M1812 229 1 6 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=52780 $D=0
M1813 230 1 6 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=57410 $D=0
M1814 231 1 6 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=62040 $D=0
M1815 232 1 6 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=66670 $D=0
M1816 7 221 229 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=52780 $D=0
M1817 7 222 230 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=57410 $D=0
M1818 7 223 231 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=62040 $D=0
M1819 7 224 232 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=66670 $D=0
M1820 233 1 8 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=52780 $D=0
M1821 234 1 9 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=57410 $D=0
M1822 235 1 10 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=62040 $D=0
M1823 236 1 11 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=66670 $D=0
M1824 8 221 233 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=52780 $D=0
M1825 9 222 234 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=57410 $D=0
M1826 10 223 235 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=62040 $D=0
M1827 11 224 236 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=66670 $D=0
M1828 241 12 233 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=52780 $D=0
M1829 242 12 234 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=57410 $D=0
M1830 243 12 235 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=62040 $D=0
M1831 244 12 236 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=66670 $D=0
M1832 237 12 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=52780 $D=0
M1833 238 12 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=57410 $D=0
M1834 239 12 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=62040 $D=0
M1835 240 12 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=66670 $D=0
M1836 245 12 229 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=52780 $D=0
M1837 246 12 230 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=57410 $D=0
M1838 247 12 231 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=62040 $D=0
M1839 248 12 232 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=66670 $D=0
M1840 225 237 245 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=52780 $D=0
M1841 226 238 246 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=57410 $D=0
M1842 227 239 247 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=62040 $D=0
M1843 228 240 248 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=66670 $D=0
M1844 249 13 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=52780 $D=0
M1845 250 13 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=57410 $D=0
M1846 251 13 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=62040 $D=0
M1847 252 13 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=66670 $D=0
M1848 253 13 245 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=52780 $D=0
M1849 254 13 246 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=57410 $D=0
M1850 255 13 247 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=62040 $D=0
M1851 256 13 248 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=66670 $D=0
M1852 241 249 253 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=52780 $D=0
M1853 242 250 254 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=57410 $D=0
M1854 243 251 255 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=62040 $D=0
M1855 244 252 256 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=66670 $D=0
M1856 257 14 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=52780 $D=0
M1857 258 14 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=57410 $D=0
M1858 259 14 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=62040 $D=0
M1859 260 14 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=66670 $D=0
M1860 261 14 8 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=52780 $D=0
M1861 262 14 9 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=57410 $D=0
M1862 263 14 10 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=62040 $D=0
M1863 264 14 11 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=66670 $D=0
M1864 15 257 261 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=52780 $D=0
M1865 16 258 262 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=57410 $D=0
M1866 17 259 263 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=62040 $D=0
M1867 18 260 264 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=66670 $D=0
M1868 265 14 19 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=52780 $D=0
M1869 266 14 20 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=57410 $D=0
M1870 267 14 21 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=62040 $D=0
M1871 268 14 22 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=66670 $D=0
M1872 269 257 265 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=52780 $D=0
M1873 270 258 266 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=57410 $D=0
M1874 271 259 267 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=62040 $D=0
M1875 272 260 268 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=66670 $D=0
M1876 277 14 273 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=52780 $D=0
M1877 278 14 274 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=57410 $D=0
M1878 279 14 275 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=62040 $D=0
M1879 280 14 276 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=66670 $D=0
M1880 253 257 277 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=52780 $D=0
M1881 254 258 278 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=57410 $D=0
M1882 255 259 279 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=62040 $D=0
M1883 256 260 280 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=66670 $D=0
M1884 285 23 277 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=52780 $D=0
M1885 286 23 278 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=57410 $D=0
M1886 287 23 279 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=62040 $D=0
M1887 288 23 280 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=66670 $D=0
M1888 281 23 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=52780 $D=0
M1889 282 23 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=57410 $D=0
M1890 283 23 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=62040 $D=0
M1891 284 23 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=66670 $D=0
M1892 289 23 265 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=52780 $D=0
M1893 290 23 266 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=57410 $D=0
M1894 291 23 267 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=62040 $D=0
M1895 292 23 268 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=66670 $D=0
M1896 261 281 289 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=52780 $D=0
M1897 262 282 290 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=57410 $D=0
M1898 263 283 291 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=62040 $D=0
M1899 264 284 292 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=66670 $D=0
M1900 293 24 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=52780 $D=0
M1901 294 24 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=57410 $D=0
M1902 295 24 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=62040 $D=0
M1903 296 24 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=66670 $D=0
M1904 297 24 289 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=52780 $D=0
M1905 298 24 290 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=57410 $D=0
M1906 299 24 291 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=62040 $D=0
M1907 300 24 292 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=66670 $D=0
M1908 285 293 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=52780 $D=0
M1909 286 294 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=57410 $D=0
M1910 287 295 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=62040 $D=0
M1911 288 296 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=66670 $D=0
M1912 191 25 301 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=52780 $D=0
M1913 192 25 302 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=57410 $D=0
M1914 193 25 303 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=62040 $D=0
M1915 194 25 304 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=66670 $D=0
M1916 305 26 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=52780 $D=0
M1917 306 26 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=57410 $D=0
M1918 307 26 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=62040 $D=0
M1919 308 26 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=66670 $D=0
M1920 309 301 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=52780 $D=0
M1921 310 302 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=57410 $D=0
M1922 311 303 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=62040 $D=0
M1923 312 304 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=66670 $D=0
M1924 191 309 1249 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=52780 $D=0
M1925 192 310 1250 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=57410 $D=0
M1926 193 311 1251 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=62040 $D=0
M1927 194 312 1252 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=66670 $D=0
M1928 313 1249 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=52780 $D=0
M1929 314 1250 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=57410 $D=0
M1930 315 1251 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=62040 $D=0
M1931 316 1252 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=66670 $D=0
M1932 309 25 313 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=52780 $D=0
M1933 310 25 314 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=57410 $D=0
M1934 311 25 315 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=62040 $D=0
M1935 312 25 316 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=66670 $D=0
M1936 313 305 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=52780 $D=0
M1937 314 306 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=57410 $D=0
M1938 315 307 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=62040 $D=0
M1939 316 308 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=66670 $D=0
M1940 325 321 313 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=52780 $D=0
M1941 326 322 314 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=57410 $D=0
M1942 327 323 315 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=62040 $D=0
M1943 328 324 316 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=66670 $D=0
M1944 321 27 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=52780 $D=0
M1945 322 27 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=57410 $D=0
M1946 323 27 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=62040 $D=0
M1947 324 27 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=66670 $D=0
M1948 191 28 329 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=52780 $D=0
M1949 192 28 330 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=57410 $D=0
M1950 193 28 331 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=62040 $D=0
M1951 194 28 332 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=66670 $D=0
M1952 333 29 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=52780 $D=0
M1953 334 29 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=57410 $D=0
M1954 335 29 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=62040 $D=0
M1955 336 29 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=66670 $D=0
M1956 337 329 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=52780 $D=0
M1957 338 330 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=57410 $D=0
M1958 339 331 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=62040 $D=0
M1959 340 332 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=66670 $D=0
M1960 191 337 1253 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=52780 $D=0
M1961 192 338 1254 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=57410 $D=0
M1962 193 339 1255 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=62040 $D=0
M1963 194 340 1256 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=66670 $D=0
M1964 341 1253 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=52780 $D=0
M1965 342 1254 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=57410 $D=0
M1966 343 1255 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=62040 $D=0
M1967 344 1256 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=66670 $D=0
M1968 337 28 341 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=52780 $D=0
M1969 338 28 342 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=57410 $D=0
M1970 339 28 343 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=62040 $D=0
M1971 340 28 344 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=66670 $D=0
M1972 341 333 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=52780 $D=0
M1973 342 334 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=57410 $D=0
M1974 343 335 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=62040 $D=0
M1975 344 336 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=66670 $D=0
M1976 325 345 341 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=52780 $D=0
M1977 326 346 342 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=57410 $D=0
M1978 327 347 343 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=62040 $D=0
M1979 328 348 344 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=66670 $D=0
M1980 345 30 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=52780 $D=0
M1981 346 30 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=57410 $D=0
M1982 347 30 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=62040 $D=0
M1983 348 30 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=66670 $D=0
M1984 191 31 349 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=52780 $D=0
M1985 192 31 350 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=57410 $D=0
M1986 193 31 351 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=62040 $D=0
M1987 194 31 352 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=66670 $D=0
M1988 353 32 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=52780 $D=0
M1989 354 32 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=57410 $D=0
M1990 355 32 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=62040 $D=0
M1991 356 32 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=66670 $D=0
M1992 357 349 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=52780 $D=0
M1993 358 350 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=57410 $D=0
M1994 359 351 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=62040 $D=0
M1995 360 352 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=66670 $D=0
M1996 191 357 1257 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=52780 $D=0
M1997 192 358 1258 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=57410 $D=0
M1998 193 359 1259 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=62040 $D=0
M1999 194 360 1260 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=66670 $D=0
M2000 361 1257 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=52780 $D=0
M2001 362 1258 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=57410 $D=0
M2002 363 1259 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=62040 $D=0
M2003 364 1260 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=66670 $D=0
M2004 357 31 361 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=52780 $D=0
M2005 358 31 362 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=57410 $D=0
M2006 359 31 363 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=62040 $D=0
M2007 360 31 364 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=66670 $D=0
M2008 361 353 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=52780 $D=0
M2009 362 354 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=57410 $D=0
M2010 363 355 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=62040 $D=0
M2011 364 356 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=66670 $D=0
M2012 325 365 361 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=52780 $D=0
M2013 326 366 362 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=57410 $D=0
M2014 327 367 363 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=62040 $D=0
M2015 328 368 364 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=66670 $D=0
M2016 365 33 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=52780 $D=0
M2017 366 33 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=57410 $D=0
M2018 367 33 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=62040 $D=0
M2019 368 33 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=66670 $D=0
M2020 191 34 369 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=52780 $D=0
M2021 192 34 370 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=57410 $D=0
M2022 193 34 371 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=62040 $D=0
M2023 194 34 372 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=66670 $D=0
M2024 373 35 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=52780 $D=0
M2025 374 35 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=57410 $D=0
M2026 375 35 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=62040 $D=0
M2027 376 35 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=66670 $D=0
M2028 377 369 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=52780 $D=0
M2029 378 370 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=57410 $D=0
M2030 379 371 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=62040 $D=0
M2031 380 372 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=66670 $D=0
M2032 191 377 1261 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=52780 $D=0
M2033 192 378 1262 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=57410 $D=0
M2034 193 379 1263 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=62040 $D=0
M2035 194 380 1264 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=66670 $D=0
M2036 381 1261 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=52780 $D=0
M2037 382 1262 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=57410 $D=0
M2038 383 1263 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=62040 $D=0
M2039 384 1264 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=66670 $D=0
M2040 377 34 381 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=52780 $D=0
M2041 378 34 382 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=57410 $D=0
M2042 379 34 383 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=62040 $D=0
M2043 380 34 384 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=66670 $D=0
M2044 381 373 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=52780 $D=0
M2045 382 374 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=57410 $D=0
M2046 383 375 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=62040 $D=0
M2047 384 376 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=66670 $D=0
M2048 325 385 381 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=52780 $D=0
M2049 326 386 382 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=57410 $D=0
M2050 327 387 383 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=62040 $D=0
M2051 328 388 384 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=66670 $D=0
M2052 385 36 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=52780 $D=0
M2053 386 36 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=57410 $D=0
M2054 387 36 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=62040 $D=0
M2055 388 36 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=66670 $D=0
M2056 191 37 389 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=52780 $D=0
M2057 192 37 390 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=57410 $D=0
M2058 193 37 391 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=62040 $D=0
M2059 194 37 392 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=66670 $D=0
M2060 393 38 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=52780 $D=0
M2061 394 38 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=57410 $D=0
M2062 395 38 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=62040 $D=0
M2063 396 38 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=66670 $D=0
M2064 397 389 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=52780 $D=0
M2065 398 390 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=57410 $D=0
M2066 399 391 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=62040 $D=0
M2067 400 392 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=66670 $D=0
M2068 191 397 1265 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=52780 $D=0
M2069 192 398 1266 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=57410 $D=0
M2070 193 399 1267 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=62040 $D=0
M2071 194 400 1268 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=66670 $D=0
M2072 401 1265 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=52780 $D=0
M2073 402 1266 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=57410 $D=0
M2074 403 1267 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=62040 $D=0
M2075 404 1268 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=66670 $D=0
M2076 397 37 401 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=52780 $D=0
M2077 398 37 402 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=57410 $D=0
M2078 399 37 403 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=62040 $D=0
M2079 400 37 404 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=66670 $D=0
M2080 401 393 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=52780 $D=0
M2081 402 394 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=57410 $D=0
M2082 403 395 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=62040 $D=0
M2083 404 396 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=66670 $D=0
M2084 325 405 401 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=52780 $D=0
M2085 326 406 402 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=57410 $D=0
M2086 327 407 403 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=62040 $D=0
M2087 328 408 404 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=66670 $D=0
M2088 405 39 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=52780 $D=0
M2089 406 39 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=57410 $D=0
M2090 407 39 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=62040 $D=0
M2091 408 39 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=66670 $D=0
M2092 191 40 409 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=52780 $D=0
M2093 192 40 410 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=57410 $D=0
M2094 193 40 411 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=62040 $D=0
M2095 194 40 412 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=66670 $D=0
M2096 413 41 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=52780 $D=0
M2097 414 41 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=57410 $D=0
M2098 415 41 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=62040 $D=0
M2099 416 41 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=66670 $D=0
M2100 417 409 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=52780 $D=0
M2101 418 410 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=57410 $D=0
M2102 419 411 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=62040 $D=0
M2103 420 412 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=66670 $D=0
M2104 191 417 1269 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=52780 $D=0
M2105 192 418 1270 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=57410 $D=0
M2106 193 419 1271 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=62040 $D=0
M2107 194 420 1272 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=66670 $D=0
M2108 421 1269 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=52780 $D=0
M2109 422 1270 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=57410 $D=0
M2110 423 1271 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=62040 $D=0
M2111 424 1272 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=66670 $D=0
M2112 417 40 421 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=52780 $D=0
M2113 418 40 422 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=57410 $D=0
M2114 419 40 423 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=62040 $D=0
M2115 420 40 424 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=66670 $D=0
M2116 421 413 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=52780 $D=0
M2117 422 414 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=57410 $D=0
M2118 423 415 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=62040 $D=0
M2119 424 416 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=66670 $D=0
M2120 325 425 421 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=52780 $D=0
M2121 326 426 422 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=57410 $D=0
M2122 327 427 423 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=62040 $D=0
M2123 328 428 424 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=66670 $D=0
M2124 425 42 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=52780 $D=0
M2125 426 42 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=57410 $D=0
M2126 427 42 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=62040 $D=0
M2127 428 42 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=66670 $D=0
M2128 191 43 429 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=52780 $D=0
M2129 192 43 430 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=57410 $D=0
M2130 193 43 431 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=62040 $D=0
M2131 194 43 432 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=66670 $D=0
M2132 433 44 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=52780 $D=0
M2133 434 44 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=57410 $D=0
M2134 435 44 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=62040 $D=0
M2135 436 44 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=66670 $D=0
M2136 437 429 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=52780 $D=0
M2137 438 430 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=57410 $D=0
M2138 439 431 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=62040 $D=0
M2139 440 432 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=66670 $D=0
M2140 191 437 1273 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=52780 $D=0
M2141 192 438 1274 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=57410 $D=0
M2142 193 439 1275 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=62040 $D=0
M2143 194 440 1276 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=66670 $D=0
M2144 441 1273 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=52780 $D=0
M2145 442 1274 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=57410 $D=0
M2146 443 1275 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=62040 $D=0
M2147 444 1276 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=66670 $D=0
M2148 437 43 441 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=52780 $D=0
M2149 438 43 442 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=57410 $D=0
M2150 439 43 443 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=62040 $D=0
M2151 440 43 444 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=66670 $D=0
M2152 441 433 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=52780 $D=0
M2153 442 434 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=57410 $D=0
M2154 443 435 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=62040 $D=0
M2155 444 436 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=66670 $D=0
M2156 325 445 441 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=52780 $D=0
M2157 326 446 442 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=57410 $D=0
M2158 327 447 443 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=62040 $D=0
M2159 328 448 444 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=66670 $D=0
M2160 445 45 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=52780 $D=0
M2161 446 45 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=57410 $D=0
M2162 447 45 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=62040 $D=0
M2163 448 45 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=66670 $D=0
M2164 191 46 449 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=52780 $D=0
M2165 192 46 450 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=57410 $D=0
M2166 193 46 451 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=62040 $D=0
M2167 194 46 452 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=66670 $D=0
M2168 453 47 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=52780 $D=0
M2169 454 47 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=57410 $D=0
M2170 455 47 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=62040 $D=0
M2171 456 47 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=66670 $D=0
M2172 457 449 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=52780 $D=0
M2173 458 450 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=57410 $D=0
M2174 459 451 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=62040 $D=0
M2175 460 452 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=66670 $D=0
M2176 191 457 1277 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=52780 $D=0
M2177 192 458 1278 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=57410 $D=0
M2178 193 459 1279 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=62040 $D=0
M2179 194 460 1280 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=66670 $D=0
M2180 461 1277 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=52780 $D=0
M2181 462 1278 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=57410 $D=0
M2182 463 1279 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=62040 $D=0
M2183 464 1280 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=66670 $D=0
M2184 457 46 461 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=52780 $D=0
M2185 458 46 462 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=57410 $D=0
M2186 459 46 463 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=62040 $D=0
M2187 460 46 464 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=66670 $D=0
M2188 461 453 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=52780 $D=0
M2189 462 454 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=57410 $D=0
M2190 463 455 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=62040 $D=0
M2191 464 456 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=66670 $D=0
M2192 325 465 461 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=52780 $D=0
M2193 326 466 462 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=57410 $D=0
M2194 327 467 463 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=62040 $D=0
M2195 328 468 464 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=66670 $D=0
M2196 465 48 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=52780 $D=0
M2197 466 48 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=57410 $D=0
M2198 467 48 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=62040 $D=0
M2199 468 48 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=66670 $D=0
M2200 191 49 469 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=52780 $D=0
M2201 192 49 470 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=57410 $D=0
M2202 193 49 471 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=62040 $D=0
M2203 194 49 472 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=66670 $D=0
M2204 473 50 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=52780 $D=0
M2205 474 50 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=57410 $D=0
M2206 475 50 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=62040 $D=0
M2207 476 50 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=66670 $D=0
M2208 477 469 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=52780 $D=0
M2209 478 470 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=57410 $D=0
M2210 479 471 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=62040 $D=0
M2211 480 472 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=66670 $D=0
M2212 191 477 1281 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=52780 $D=0
M2213 192 478 1282 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=57410 $D=0
M2214 193 479 1283 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=62040 $D=0
M2215 194 480 1284 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=66670 $D=0
M2216 481 1281 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=52780 $D=0
M2217 482 1282 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=57410 $D=0
M2218 483 1283 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=62040 $D=0
M2219 484 1284 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=66670 $D=0
M2220 477 49 481 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=52780 $D=0
M2221 478 49 482 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=57410 $D=0
M2222 479 49 483 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=62040 $D=0
M2223 480 49 484 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=66670 $D=0
M2224 481 473 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=52780 $D=0
M2225 482 474 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=57410 $D=0
M2226 483 475 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=62040 $D=0
M2227 484 476 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=66670 $D=0
M2228 325 485 481 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=52780 $D=0
M2229 326 486 482 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=57410 $D=0
M2230 327 487 483 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=62040 $D=0
M2231 328 488 484 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=66670 $D=0
M2232 485 51 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=52780 $D=0
M2233 486 51 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=57410 $D=0
M2234 487 51 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=62040 $D=0
M2235 488 51 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=66670 $D=0
M2236 191 52 489 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=52780 $D=0
M2237 192 52 490 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=57410 $D=0
M2238 193 52 491 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=62040 $D=0
M2239 194 52 492 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=66670 $D=0
M2240 493 53 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=52780 $D=0
M2241 494 53 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=57410 $D=0
M2242 495 53 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=62040 $D=0
M2243 496 53 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=66670 $D=0
M2244 497 489 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=52780 $D=0
M2245 498 490 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=57410 $D=0
M2246 499 491 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=62040 $D=0
M2247 500 492 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=66670 $D=0
M2248 191 497 1285 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=52780 $D=0
M2249 192 498 1286 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=57410 $D=0
M2250 193 499 1287 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=62040 $D=0
M2251 194 500 1288 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=66670 $D=0
M2252 501 1285 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=52780 $D=0
M2253 502 1286 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=57410 $D=0
M2254 503 1287 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=62040 $D=0
M2255 504 1288 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=66670 $D=0
M2256 497 52 501 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=52780 $D=0
M2257 498 52 502 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=57410 $D=0
M2258 499 52 503 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=62040 $D=0
M2259 500 52 504 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=66670 $D=0
M2260 501 493 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=52780 $D=0
M2261 502 494 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=57410 $D=0
M2262 503 495 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=62040 $D=0
M2263 504 496 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=66670 $D=0
M2264 325 505 501 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=52780 $D=0
M2265 326 506 502 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=57410 $D=0
M2266 327 507 503 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=62040 $D=0
M2267 328 508 504 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=66670 $D=0
M2268 505 54 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=52780 $D=0
M2269 506 54 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=57410 $D=0
M2270 507 54 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=62040 $D=0
M2271 508 54 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=66670 $D=0
M2272 191 55 509 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=52780 $D=0
M2273 192 55 510 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=57410 $D=0
M2274 193 55 511 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=62040 $D=0
M2275 194 55 512 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=66670 $D=0
M2276 513 56 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=52780 $D=0
M2277 514 56 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=57410 $D=0
M2278 515 56 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=62040 $D=0
M2279 516 56 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=66670 $D=0
M2280 517 509 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=52780 $D=0
M2281 518 510 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=57410 $D=0
M2282 519 511 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=62040 $D=0
M2283 520 512 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=66670 $D=0
M2284 191 517 1289 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=52780 $D=0
M2285 192 518 1290 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=57410 $D=0
M2286 193 519 1291 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=62040 $D=0
M2287 194 520 1292 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=66670 $D=0
M2288 521 1289 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=52780 $D=0
M2289 522 1290 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=57410 $D=0
M2290 523 1291 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=62040 $D=0
M2291 524 1292 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=66670 $D=0
M2292 517 55 521 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=52780 $D=0
M2293 518 55 522 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=57410 $D=0
M2294 519 55 523 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=62040 $D=0
M2295 520 55 524 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=66670 $D=0
M2296 521 513 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=52780 $D=0
M2297 522 514 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=57410 $D=0
M2298 523 515 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=62040 $D=0
M2299 524 516 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=66670 $D=0
M2300 325 525 521 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=52780 $D=0
M2301 326 526 522 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=57410 $D=0
M2302 327 527 523 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=62040 $D=0
M2303 328 528 524 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=66670 $D=0
M2304 525 57 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=52780 $D=0
M2305 526 57 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=57410 $D=0
M2306 527 57 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=62040 $D=0
M2307 528 57 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=66670 $D=0
M2308 191 58 529 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=52780 $D=0
M2309 192 58 530 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=57410 $D=0
M2310 193 58 531 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=62040 $D=0
M2311 194 58 532 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=66670 $D=0
M2312 533 59 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=52780 $D=0
M2313 534 59 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=57410 $D=0
M2314 535 59 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=62040 $D=0
M2315 536 59 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=66670 $D=0
M2316 537 529 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=52780 $D=0
M2317 538 530 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=57410 $D=0
M2318 539 531 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=62040 $D=0
M2319 540 532 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=66670 $D=0
M2320 191 537 1293 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=52780 $D=0
M2321 192 538 1294 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=57410 $D=0
M2322 193 539 1295 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=62040 $D=0
M2323 194 540 1296 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=66670 $D=0
M2324 541 1293 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=52780 $D=0
M2325 542 1294 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=57410 $D=0
M2326 543 1295 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=62040 $D=0
M2327 544 1296 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=66670 $D=0
M2328 537 58 541 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=52780 $D=0
M2329 538 58 542 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=57410 $D=0
M2330 539 58 543 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=62040 $D=0
M2331 540 58 544 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=66670 $D=0
M2332 541 533 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=52780 $D=0
M2333 542 534 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=57410 $D=0
M2334 543 535 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=62040 $D=0
M2335 544 536 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=66670 $D=0
M2336 325 545 541 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=52780 $D=0
M2337 326 546 542 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=57410 $D=0
M2338 327 547 543 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=62040 $D=0
M2339 328 548 544 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=66670 $D=0
M2340 545 60 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=52780 $D=0
M2341 546 60 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=57410 $D=0
M2342 547 60 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=62040 $D=0
M2343 548 60 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=66670 $D=0
M2344 191 61 549 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=52780 $D=0
M2345 192 61 550 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=57410 $D=0
M2346 193 61 551 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=62040 $D=0
M2347 194 61 552 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=66670 $D=0
M2348 553 62 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=52780 $D=0
M2349 554 62 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=57410 $D=0
M2350 555 62 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=62040 $D=0
M2351 556 62 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=66670 $D=0
M2352 557 549 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=52780 $D=0
M2353 558 550 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=57410 $D=0
M2354 559 551 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=62040 $D=0
M2355 560 552 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=66670 $D=0
M2356 191 557 1297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=52780 $D=0
M2357 192 558 1298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=57410 $D=0
M2358 193 559 1299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=62040 $D=0
M2359 194 560 1300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=66670 $D=0
M2360 561 1297 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=52780 $D=0
M2361 562 1298 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=57410 $D=0
M2362 563 1299 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=62040 $D=0
M2363 564 1300 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=66670 $D=0
M2364 557 61 561 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=52780 $D=0
M2365 558 61 562 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=57410 $D=0
M2366 559 61 563 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=62040 $D=0
M2367 560 61 564 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=66670 $D=0
M2368 561 553 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=52780 $D=0
M2369 562 554 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=57410 $D=0
M2370 563 555 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=62040 $D=0
M2371 564 556 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=66670 $D=0
M2372 325 565 561 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=52780 $D=0
M2373 326 566 562 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=57410 $D=0
M2374 327 567 563 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=62040 $D=0
M2375 328 568 564 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=66670 $D=0
M2376 565 63 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=52780 $D=0
M2377 566 63 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=57410 $D=0
M2378 567 63 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=62040 $D=0
M2379 568 63 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=66670 $D=0
M2380 191 64 569 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=52780 $D=0
M2381 192 64 570 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=57410 $D=0
M2382 193 64 571 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=62040 $D=0
M2383 194 64 572 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=66670 $D=0
M2384 573 65 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=52780 $D=0
M2385 574 65 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=57410 $D=0
M2386 575 65 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=62040 $D=0
M2387 576 65 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=66670 $D=0
M2388 577 569 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=52780 $D=0
M2389 578 570 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=57410 $D=0
M2390 579 571 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=62040 $D=0
M2391 580 572 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=66670 $D=0
M2392 191 577 1301 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=52780 $D=0
M2393 192 578 1302 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=57410 $D=0
M2394 193 579 1303 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=62040 $D=0
M2395 194 580 1304 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=66670 $D=0
M2396 581 1301 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=52780 $D=0
M2397 582 1302 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=57410 $D=0
M2398 583 1303 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=62040 $D=0
M2399 584 1304 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=66670 $D=0
M2400 577 64 581 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=52780 $D=0
M2401 578 64 582 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=57410 $D=0
M2402 579 64 583 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=62040 $D=0
M2403 580 64 584 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=66670 $D=0
M2404 581 573 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=52780 $D=0
M2405 582 574 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=57410 $D=0
M2406 583 575 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=62040 $D=0
M2407 584 576 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=66670 $D=0
M2408 325 585 581 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=52780 $D=0
M2409 326 586 582 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=57410 $D=0
M2410 327 587 583 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=62040 $D=0
M2411 328 588 584 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=66670 $D=0
M2412 585 66 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=52780 $D=0
M2413 586 66 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=57410 $D=0
M2414 587 66 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=62040 $D=0
M2415 588 66 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=66670 $D=0
M2416 191 67 589 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=52780 $D=0
M2417 192 67 590 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=57410 $D=0
M2418 193 67 591 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=62040 $D=0
M2419 194 67 592 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=66670 $D=0
M2420 593 68 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=52780 $D=0
M2421 594 68 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=57410 $D=0
M2422 595 68 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=62040 $D=0
M2423 596 68 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=66670 $D=0
M2424 597 589 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=52780 $D=0
M2425 598 590 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=57410 $D=0
M2426 599 591 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=62040 $D=0
M2427 600 592 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=66670 $D=0
M2428 191 597 1305 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=52780 $D=0
M2429 192 598 1306 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=57410 $D=0
M2430 193 599 1307 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=62040 $D=0
M2431 194 600 1308 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=66670 $D=0
M2432 601 1305 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=52780 $D=0
M2433 602 1306 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=57410 $D=0
M2434 603 1307 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=62040 $D=0
M2435 604 1308 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=66670 $D=0
M2436 597 67 601 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=52780 $D=0
M2437 598 67 602 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=57410 $D=0
M2438 599 67 603 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=62040 $D=0
M2439 600 67 604 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=66670 $D=0
M2440 601 593 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=52780 $D=0
M2441 602 594 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=57410 $D=0
M2442 603 595 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=62040 $D=0
M2443 604 596 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=66670 $D=0
M2444 325 605 601 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=52780 $D=0
M2445 326 606 602 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=57410 $D=0
M2446 327 607 603 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=62040 $D=0
M2447 328 608 604 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=66670 $D=0
M2448 605 69 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=52780 $D=0
M2449 606 69 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=57410 $D=0
M2450 607 69 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=62040 $D=0
M2451 608 69 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=66670 $D=0
M2452 191 70 609 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=52780 $D=0
M2453 192 70 610 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=57410 $D=0
M2454 193 70 611 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=62040 $D=0
M2455 194 70 612 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=66670 $D=0
M2456 613 71 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=52780 $D=0
M2457 614 71 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=57410 $D=0
M2458 615 71 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=62040 $D=0
M2459 616 71 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=66670 $D=0
M2460 617 609 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=52780 $D=0
M2461 618 610 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=57410 $D=0
M2462 619 611 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=62040 $D=0
M2463 620 612 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=66670 $D=0
M2464 191 617 1309 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=52780 $D=0
M2465 192 618 1310 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=57410 $D=0
M2466 193 619 1311 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=62040 $D=0
M2467 194 620 1312 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=66670 $D=0
M2468 621 1309 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=52780 $D=0
M2469 622 1310 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=57410 $D=0
M2470 623 1311 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=62040 $D=0
M2471 624 1312 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=66670 $D=0
M2472 617 70 621 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=52780 $D=0
M2473 618 70 622 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=57410 $D=0
M2474 619 70 623 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=62040 $D=0
M2475 620 70 624 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=66670 $D=0
M2476 621 613 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=52780 $D=0
M2477 622 614 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=57410 $D=0
M2478 623 615 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=62040 $D=0
M2479 624 616 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=66670 $D=0
M2480 325 625 621 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=52780 $D=0
M2481 326 626 622 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=57410 $D=0
M2482 327 627 623 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=62040 $D=0
M2483 328 628 624 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=66670 $D=0
M2484 625 72 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=52780 $D=0
M2485 626 72 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=57410 $D=0
M2486 627 72 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=62040 $D=0
M2487 628 72 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=66670 $D=0
M2488 191 73 629 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=52780 $D=0
M2489 192 73 630 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=57410 $D=0
M2490 193 73 631 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=62040 $D=0
M2491 194 73 632 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=66670 $D=0
M2492 633 74 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=52780 $D=0
M2493 634 74 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=57410 $D=0
M2494 635 74 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=62040 $D=0
M2495 636 74 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=66670 $D=0
M2496 637 629 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=52780 $D=0
M2497 638 630 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=57410 $D=0
M2498 639 631 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=62040 $D=0
M2499 640 632 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=66670 $D=0
M2500 191 637 1313 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=52780 $D=0
M2501 192 638 1314 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=57410 $D=0
M2502 193 639 1315 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=62040 $D=0
M2503 194 640 1316 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=66670 $D=0
M2504 641 1313 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=52780 $D=0
M2505 642 1314 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=57410 $D=0
M2506 643 1315 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=62040 $D=0
M2507 644 1316 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=66670 $D=0
M2508 637 73 641 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=52780 $D=0
M2509 638 73 642 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=57410 $D=0
M2510 639 73 643 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=62040 $D=0
M2511 640 73 644 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=66670 $D=0
M2512 641 633 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=52780 $D=0
M2513 642 634 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=57410 $D=0
M2514 643 635 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=62040 $D=0
M2515 644 636 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=66670 $D=0
M2516 325 645 641 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=52780 $D=0
M2517 326 646 642 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=57410 $D=0
M2518 327 647 643 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=62040 $D=0
M2519 328 648 644 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=66670 $D=0
M2520 645 75 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=52780 $D=0
M2521 646 75 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=57410 $D=0
M2522 647 75 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=62040 $D=0
M2523 648 75 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=66670 $D=0
M2524 191 76 649 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=52780 $D=0
M2525 192 76 650 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=57410 $D=0
M2526 193 76 651 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=62040 $D=0
M2527 194 76 652 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=66670 $D=0
M2528 653 77 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=52780 $D=0
M2529 654 77 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=57410 $D=0
M2530 655 77 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=62040 $D=0
M2531 656 77 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=66670 $D=0
M2532 657 649 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=52780 $D=0
M2533 658 650 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=57410 $D=0
M2534 659 651 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=62040 $D=0
M2535 660 652 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=66670 $D=0
M2536 191 657 1317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=52780 $D=0
M2537 192 658 1318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=57410 $D=0
M2538 193 659 1319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=62040 $D=0
M2539 194 660 1320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=66670 $D=0
M2540 661 1317 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=52780 $D=0
M2541 662 1318 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=57410 $D=0
M2542 663 1319 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=62040 $D=0
M2543 664 1320 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=66670 $D=0
M2544 657 76 661 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=52780 $D=0
M2545 658 76 662 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=57410 $D=0
M2546 659 76 663 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=62040 $D=0
M2547 660 76 664 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=66670 $D=0
M2548 661 653 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=52780 $D=0
M2549 662 654 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=57410 $D=0
M2550 663 655 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=62040 $D=0
M2551 664 656 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=66670 $D=0
M2552 325 665 661 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=52780 $D=0
M2553 326 666 662 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=57410 $D=0
M2554 327 667 663 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=62040 $D=0
M2555 328 668 664 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=66670 $D=0
M2556 665 78 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=52780 $D=0
M2557 666 78 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=57410 $D=0
M2558 667 78 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=62040 $D=0
M2559 668 78 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=66670 $D=0
M2560 191 79 669 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=52780 $D=0
M2561 192 79 670 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=57410 $D=0
M2562 193 79 671 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=62040 $D=0
M2563 194 79 672 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=66670 $D=0
M2564 673 80 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=52780 $D=0
M2565 674 80 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=57410 $D=0
M2566 675 80 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=62040 $D=0
M2567 676 80 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=66670 $D=0
M2568 677 669 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=52780 $D=0
M2569 678 670 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=57410 $D=0
M2570 679 671 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=62040 $D=0
M2571 680 672 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=66670 $D=0
M2572 191 677 1321 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=52780 $D=0
M2573 192 678 1322 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=57410 $D=0
M2574 193 679 1323 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=62040 $D=0
M2575 194 680 1324 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=66670 $D=0
M2576 681 1321 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=52780 $D=0
M2577 682 1322 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=57410 $D=0
M2578 683 1323 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=62040 $D=0
M2579 684 1324 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=66670 $D=0
M2580 677 79 681 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=52780 $D=0
M2581 678 79 682 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=57410 $D=0
M2582 679 79 683 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=62040 $D=0
M2583 680 79 684 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=66670 $D=0
M2584 681 673 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=52780 $D=0
M2585 682 674 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=57410 $D=0
M2586 683 675 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=62040 $D=0
M2587 684 676 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=66670 $D=0
M2588 325 685 681 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=52780 $D=0
M2589 326 686 682 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=57410 $D=0
M2590 327 687 683 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=62040 $D=0
M2591 328 688 684 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=66670 $D=0
M2592 685 81 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=52780 $D=0
M2593 686 81 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=57410 $D=0
M2594 687 81 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=62040 $D=0
M2595 688 81 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=66670 $D=0
M2596 191 82 689 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=52780 $D=0
M2597 192 82 690 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=57410 $D=0
M2598 193 82 691 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=62040 $D=0
M2599 194 82 692 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=66670 $D=0
M2600 693 83 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=52780 $D=0
M2601 694 83 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=57410 $D=0
M2602 695 83 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=62040 $D=0
M2603 696 83 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=66670 $D=0
M2604 697 689 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=52780 $D=0
M2605 698 690 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=57410 $D=0
M2606 699 691 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=62040 $D=0
M2607 700 692 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=66670 $D=0
M2608 191 697 1325 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=52780 $D=0
M2609 192 698 1326 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=57410 $D=0
M2610 193 699 1327 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=62040 $D=0
M2611 194 700 1328 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=66670 $D=0
M2612 701 1325 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=52780 $D=0
M2613 702 1326 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=57410 $D=0
M2614 703 1327 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=62040 $D=0
M2615 704 1328 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=66670 $D=0
M2616 697 82 701 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=52780 $D=0
M2617 698 82 702 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=57410 $D=0
M2618 699 82 703 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=62040 $D=0
M2619 700 82 704 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=66670 $D=0
M2620 701 693 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=52780 $D=0
M2621 702 694 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=57410 $D=0
M2622 703 695 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=62040 $D=0
M2623 704 696 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=66670 $D=0
M2624 325 705 701 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=52780 $D=0
M2625 326 706 702 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=57410 $D=0
M2626 327 707 703 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=62040 $D=0
M2627 328 708 704 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=66670 $D=0
M2628 705 84 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=52780 $D=0
M2629 706 84 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=57410 $D=0
M2630 707 84 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=62040 $D=0
M2631 708 84 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=66670 $D=0
M2632 191 85 709 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=52780 $D=0
M2633 192 85 710 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=57410 $D=0
M2634 193 85 711 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=62040 $D=0
M2635 194 85 712 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=66670 $D=0
M2636 713 86 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=52780 $D=0
M2637 714 86 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=57410 $D=0
M2638 715 86 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=62040 $D=0
M2639 716 86 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=66670 $D=0
M2640 717 709 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=52780 $D=0
M2641 718 710 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=57410 $D=0
M2642 719 711 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=62040 $D=0
M2643 720 712 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=66670 $D=0
M2644 191 717 1329 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=52780 $D=0
M2645 192 718 1330 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=57410 $D=0
M2646 193 719 1331 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=62040 $D=0
M2647 194 720 1332 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=66670 $D=0
M2648 721 1329 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=52780 $D=0
M2649 722 1330 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=57410 $D=0
M2650 723 1331 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=62040 $D=0
M2651 724 1332 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=66670 $D=0
M2652 717 85 721 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=52780 $D=0
M2653 718 85 722 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=57410 $D=0
M2654 719 85 723 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=62040 $D=0
M2655 720 85 724 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=66670 $D=0
M2656 721 713 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=52780 $D=0
M2657 722 714 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=57410 $D=0
M2658 723 715 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=62040 $D=0
M2659 724 716 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=66670 $D=0
M2660 325 725 721 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=52780 $D=0
M2661 326 726 722 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=57410 $D=0
M2662 327 727 723 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=62040 $D=0
M2663 328 728 724 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=66670 $D=0
M2664 725 87 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=52780 $D=0
M2665 726 87 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=57410 $D=0
M2666 727 87 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=62040 $D=0
M2667 728 87 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=66670 $D=0
M2668 191 88 729 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=52780 $D=0
M2669 192 88 730 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=57410 $D=0
M2670 193 88 731 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=62040 $D=0
M2671 194 88 732 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=66670 $D=0
M2672 733 89 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=52780 $D=0
M2673 734 89 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=57410 $D=0
M2674 735 89 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=62040 $D=0
M2675 736 89 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=66670 $D=0
M2676 737 729 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=52780 $D=0
M2677 738 730 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=57410 $D=0
M2678 739 731 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=62040 $D=0
M2679 740 732 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=66670 $D=0
M2680 191 737 1333 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=52780 $D=0
M2681 192 738 1334 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=57410 $D=0
M2682 193 739 1335 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=62040 $D=0
M2683 194 740 1336 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=66670 $D=0
M2684 741 1333 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=52780 $D=0
M2685 742 1334 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=57410 $D=0
M2686 743 1335 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=62040 $D=0
M2687 744 1336 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=66670 $D=0
M2688 737 88 741 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=52780 $D=0
M2689 738 88 742 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=57410 $D=0
M2690 739 88 743 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=62040 $D=0
M2691 740 88 744 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=66670 $D=0
M2692 741 733 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=52780 $D=0
M2693 742 734 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=57410 $D=0
M2694 743 735 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=62040 $D=0
M2695 744 736 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=66670 $D=0
M2696 325 745 741 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=52780 $D=0
M2697 326 746 742 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=57410 $D=0
M2698 327 747 743 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=62040 $D=0
M2699 328 748 744 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=66670 $D=0
M2700 745 90 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=52780 $D=0
M2701 746 90 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=57410 $D=0
M2702 747 90 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=62040 $D=0
M2703 748 90 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=66670 $D=0
M2704 191 91 749 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=52780 $D=0
M2705 192 91 750 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=57410 $D=0
M2706 193 91 751 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=62040 $D=0
M2707 194 91 752 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=66670 $D=0
M2708 753 92 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=52780 $D=0
M2709 754 92 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=57410 $D=0
M2710 755 92 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=62040 $D=0
M2711 756 92 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=66670 $D=0
M2712 757 749 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=52780 $D=0
M2713 758 750 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=57410 $D=0
M2714 759 751 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=62040 $D=0
M2715 760 752 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=66670 $D=0
M2716 191 757 1337 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=52780 $D=0
M2717 192 758 1338 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=57410 $D=0
M2718 193 759 1339 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=62040 $D=0
M2719 194 760 1340 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=66670 $D=0
M2720 761 1337 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=52780 $D=0
M2721 762 1338 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=57410 $D=0
M2722 763 1339 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=62040 $D=0
M2723 764 1340 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=66670 $D=0
M2724 757 91 761 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=52780 $D=0
M2725 758 91 762 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=57410 $D=0
M2726 759 91 763 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=62040 $D=0
M2727 760 91 764 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=66670 $D=0
M2728 761 753 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=52780 $D=0
M2729 762 754 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=57410 $D=0
M2730 763 755 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=62040 $D=0
M2731 764 756 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=66670 $D=0
M2732 325 765 761 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=52780 $D=0
M2733 326 766 762 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=57410 $D=0
M2734 327 767 763 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=62040 $D=0
M2735 328 768 764 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=66670 $D=0
M2736 765 93 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=52780 $D=0
M2737 766 93 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=57410 $D=0
M2738 767 93 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=62040 $D=0
M2739 768 93 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=66670 $D=0
M2740 191 94 769 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=52780 $D=0
M2741 192 94 770 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=57410 $D=0
M2742 193 94 771 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=62040 $D=0
M2743 194 94 772 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=66670 $D=0
M2744 773 95 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=52780 $D=0
M2745 774 95 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=57410 $D=0
M2746 775 95 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=62040 $D=0
M2747 776 95 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=66670 $D=0
M2748 777 769 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=52780 $D=0
M2749 778 770 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=57410 $D=0
M2750 779 771 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=62040 $D=0
M2751 780 772 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=66670 $D=0
M2752 191 777 1341 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=52780 $D=0
M2753 192 778 1342 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=57410 $D=0
M2754 193 779 1343 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=62040 $D=0
M2755 194 780 1344 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=66670 $D=0
M2756 781 1341 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=52780 $D=0
M2757 782 1342 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=57410 $D=0
M2758 783 1343 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=62040 $D=0
M2759 784 1344 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=66670 $D=0
M2760 777 94 781 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=52780 $D=0
M2761 778 94 782 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=57410 $D=0
M2762 779 94 783 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=62040 $D=0
M2763 780 94 784 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=66670 $D=0
M2764 781 773 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=52780 $D=0
M2765 782 774 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=57410 $D=0
M2766 783 775 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=62040 $D=0
M2767 784 776 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=66670 $D=0
M2768 325 785 781 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=52780 $D=0
M2769 326 786 782 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=57410 $D=0
M2770 327 787 783 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=62040 $D=0
M2771 328 788 784 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=66670 $D=0
M2772 785 96 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=52780 $D=0
M2773 786 96 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=57410 $D=0
M2774 787 96 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=62040 $D=0
M2775 788 96 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=66670 $D=0
M2776 191 97 789 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=52780 $D=0
M2777 192 97 790 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=57410 $D=0
M2778 193 97 791 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=62040 $D=0
M2779 194 97 792 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=66670 $D=0
M2780 793 98 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=52780 $D=0
M2781 794 98 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=57410 $D=0
M2782 795 98 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=62040 $D=0
M2783 796 98 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=66670 $D=0
M2784 797 789 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=52780 $D=0
M2785 798 790 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=57410 $D=0
M2786 799 791 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=62040 $D=0
M2787 800 792 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=66670 $D=0
M2788 191 797 1345 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=52780 $D=0
M2789 192 798 1346 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=57410 $D=0
M2790 193 799 1347 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=62040 $D=0
M2791 194 800 1348 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=66670 $D=0
M2792 801 1345 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=52780 $D=0
M2793 802 1346 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=57410 $D=0
M2794 803 1347 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=62040 $D=0
M2795 804 1348 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=66670 $D=0
M2796 797 97 801 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=52780 $D=0
M2797 798 97 802 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=57410 $D=0
M2798 799 97 803 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=62040 $D=0
M2799 800 97 804 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=66670 $D=0
M2800 801 793 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=52780 $D=0
M2801 802 794 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=57410 $D=0
M2802 803 795 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=62040 $D=0
M2803 804 796 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=66670 $D=0
M2804 325 805 801 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=52780 $D=0
M2805 326 806 802 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=57410 $D=0
M2806 327 807 803 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=62040 $D=0
M2807 328 808 804 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=66670 $D=0
M2808 805 99 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=52780 $D=0
M2809 806 99 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=57410 $D=0
M2810 807 99 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=62040 $D=0
M2811 808 99 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=66670 $D=0
M2812 191 100 809 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=52780 $D=0
M2813 192 100 810 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=57410 $D=0
M2814 193 100 811 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=62040 $D=0
M2815 194 100 812 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=66670 $D=0
M2816 813 101 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=52780 $D=0
M2817 814 101 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=57410 $D=0
M2818 815 101 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=62040 $D=0
M2819 816 101 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=66670 $D=0
M2820 817 809 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=52780 $D=0
M2821 818 810 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=57410 $D=0
M2822 819 811 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=62040 $D=0
M2823 820 812 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=66670 $D=0
M2824 191 817 1349 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=52780 $D=0
M2825 192 818 1350 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=57410 $D=0
M2826 193 819 1351 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=62040 $D=0
M2827 194 820 1352 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=66670 $D=0
M2828 821 1349 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=52780 $D=0
M2829 822 1350 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=57410 $D=0
M2830 823 1351 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=62040 $D=0
M2831 824 1352 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=66670 $D=0
M2832 817 100 821 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=52780 $D=0
M2833 818 100 822 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=57410 $D=0
M2834 819 100 823 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=62040 $D=0
M2835 820 100 824 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=66670 $D=0
M2836 821 813 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=52780 $D=0
M2837 822 814 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=57410 $D=0
M2838 823 815 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=62040 $D=0
M2839 824 816 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=66670 $D=0
M2840 325 825 821 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=52780 $D=0
M2841 326 826 822 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=57410 $D=0
M2842 327 827 823 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=62040 $D=0
M2843 328 828 824 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=66670 $D=0
M2844 825 102 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=52780 $D=0
M2845 826 102 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=57410 $D=0
M2846 827 102 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=62040 $D=0
M2847 828 102 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=66670 $D=0
M2848 191 103 829 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=52780 $D=0
M2849 192 103 830 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=57410 $D=0
M2850 193 103 831 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=62040 $D=0
M2851 194 103 832 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=66670 $D=0
M2852 833 104 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=52780 $D=0
M2853 834 104 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=57410 $D=0
M2854 835 104 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=62040 $D=0
M2855 836 104 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=66670 $D=0
M2856 837 829 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=52780 $D=0
M2857 838 830 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=57410 $D=0
M2858 839 831 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=62040 $D=0
M2859 840 832 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=66670 $D=0
M2860 191 837 1353 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=52780 $D=0
M2861 192 838 1354 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=57410 $D=0
M2862 193 839 1355 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=62040 $D=0
M2863 194 840 1356 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=66670 $D=0
M2864 841 1353 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=52780 $D=0
M2865 842 1354 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=57410 $D=0
M2866 843 1355 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=62040 $D=0
M2867 844 1356 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=66670 $D=0
M2868 837 103 841 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=52780 $D=0
M2869 838 103 842 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=57410 $D=0
M2870 839 103 843 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=62040 $D=0
M2871 840 103 844 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=66670 $D=0
M2872 841 833 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=52780 $D=0
M2873 842 834 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=57410 $D=0
M2874 843 835 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=62040 $D=0
M2875 844 836 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=66670 $D=0
M2876 325 845 841 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=52780 $D=0
M2877 326 846 842 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=57410 $D=0
M2878 327 847 843 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=62040 $D=0
M2879 328 848 844 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=66670 $D=0
M2880 845 105 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=52780 $D=0
M2881 846 105 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=57410 $D=0
M2882 847 105 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=62040 $D=0
M2883 848 105 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=66670 $D=0
M2884 191 106 849 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=52780 $D=0
M2885 192 106 850 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=57410 $D=0
M2886 193 106 851 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=62040 $D=0
M2887 194 106 852 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=66670 $D=0
M2888 853 107 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=52780 $D=0
M2889 854 107 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=57410 $D=0
M2890 855 107 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=62040 $D=0
M2891 856 107 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=66670 $D=0
M2892 857 849 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=52780 $D=0
M2893 858 850 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=57410 $D=0
M2894 859 851 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=62040 $D=0
M2895 860 852 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=66670 $D=0
M2896 191 857 1357 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=52780 $D=0
M2897 192 858 1358 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=57410 $D=0
M2898 193 859 1359 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=62040 $D=0
M2899 194 860 1360 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=66670 $D=0
M2900 861 1357 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=52780 $D=0
M2901 862 1358 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=57410 $D=0
M2902 863 1359 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=62040 $D=0
M2903 864 1360 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=66670 $D=0
M2904 857 106 861 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=52780 $D=0
M2905 858 106 862 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=57410 $D=0
M2906 859 106 863 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=62040 $D=0
M2907 860 106 864 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=66670 $D=0
M2908 861 853 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=52780 $D=0
M2909 862 854 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=57410 $D=0
M2910 863 855 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=62040 $D=0
M2911 864 856 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=66670 $D=0
M2912 325 865 861 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=52780 $D=0
M2913 326 866 862 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=57410 $D=0
M2914 327 867 863 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=62040 $D=0
M2915 328 868 864 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=66670 $D=0
M2916 865 108 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=52780 $D=0
M2917 866 108 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=57410 $D=0
M2918 867 108 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=62040 $D=0
M2919 868 108 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=66670 $D=0
M2920 191 109 869 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=52780 $D=0
M2921 192 109 870 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=57410 $D=0
M2922 193 109 871 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=62040 $D=0
M2923 194 109 872 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=66670 $D=0
M2924 873 110 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=52780 $D=0
M2925 874 110 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=57410 $D=0
M2926 875 110 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=62040 $D=0
M2927 876 110 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=66670 $D=0
M2928 877 869 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=52780 $D=0
M2929 878 870 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=57410 $D=0
M2930 879 871 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=62040 $D=0
M2931 880 872 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=66670 $D=0
M2932 191 877 1361 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=52780 $D=0
M2933 192 878 1362 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=57410 $D=0
M2934 193 879 1363 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=62040 $D=0
M2935 194 880 1364 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=66670 $D=0
M2936 881 1361 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=52780 $D=0
M2937 882 1362 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=57410 $D=0
M2938 883 1363 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=62040 $D=0
M2939 884 1364 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=66670 $D=0
M2940 877 109 881 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=52780 $D=0
M2941 878 109 882 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=57410 $D=0
M2942 879 109 883 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=62040 $D=0
M2943 880 109 884 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=66670 $D=0
M2944 881 873 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=52780 $D=0
M2945 882 874 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=57410 $D=0
M2946 883 875 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=62040 $D=0
M2947 884 876 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=66670 $D=0
M2948 325 885 881 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=52780 $D=0
M2949 326 886 882 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=57410 $D=0
M2950 327 887 883 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=62040 $D=0
M2951 328 888 884 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=66670 $D=0
M2952 885 111 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=52780 $D=0
M2953 886 111 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=57410 $D=0
M2954 887 111 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=62040 $D=0
M2955 888 111 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=66670 $D=0
M2956 191 112 889 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=52780 $D=0
M2957 192 112 890 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=57410 $D=0
M2958 193 112 891 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=62040 $D=0
M2959 194 112 892 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=66670 $D=0
M2960 893 113 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=52780 $D=0
M2961 894 113 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=57410 $D=0
M2962 895 113 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=62040 $D=0
M2963 896 113 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=66670 $D=0
M2964 897 889 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=52780 $D=0
M2965 898 890 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=57410 $D=0
M2966 899 891 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=62040 $D=0
M2967 900 892 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=66670 $D=0
M2968 191 897 1365 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=52780 $D=0
M2969 192 898 1366 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=57410 $D=0
M2970 193 899 1367 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=62040 $D=0
M2971 194 900 1368 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=66670 $D=0
M2972 901 1365 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=52780 $D=0
M2973 902 1366 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=57410 $D=0
M2974 903 1367 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=62040 $D=0
M2975 904 1368 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=66670 $D=0
M2976 897 112 901 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=52780 $D=0
M2977 898 112 902 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=57410 $D=0
M2978 899 112 903 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=62040 $D=0
M2979 900 112 904 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=66670 $D=0
M2980 901 893 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=52780 $D=0
M2981 902 894 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=57410 $D=0
M2982 903 895 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=62040 $D=0
M2983 904 896 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=66670 $D=0
M2984 325 905 901 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=52780 $D=0
M2985 326 906 902 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=57410 $D=0
M2986 327 907 903 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=62040 $D=0
M2987 328 908 904 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=66670 $D=0
M2988 905 116 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=52780 $D=0
M2989 906 116 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=57410 $D=0
M2990 907 116 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=62040 $D=0
M2991 908 116 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=66670 $D=0
M2992 191 117 909 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=52780 $D=0
M2993 192 117 910 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=57410 $D=0
M2994 193 117 911 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=62040 $D=0
M2995 194 117 912 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=66670 $D=0
M2996 913 118 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=52780 $D=0
M2997 914 118 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=57410 $D=0
M2998 915 118 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=62040 $D=0
M2999 916 118 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=66670 $D=0
M3000 917 909 297 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=52780 $D=0
M3001 918 910 298 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=57410 $D=0
M3002 919 911 299 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=62040 $D=0
M3003 920 912 300 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=66670 $D=0
M3004 191 917 1369 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=52780 $D=0
M3005 192 918 1370 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=57410 $D=0
M3006 193 919 1371 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=62040 $D=0
M3007 194 920 1372 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=66670 $D=0
M3008 921 1369 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=52780 $D=0
M3009 922 1370 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=57410 $D=0
M3010 923 1371 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=62040 $D=0
M3011 924 1372 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=66670 $D=0
M3012 917 117 921 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=52780 $D=0
M3013 918 117 922 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=57410 $D=0
M3014 919 117 923 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=62040 $D=0
M3015 920 117 924 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=66670 $D=0
M3016 921 913 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=52780 $D=0
M3017 922 914 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=57410 $D=0
M3018 923 915 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=62040 $D=0
M3019 924 916 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=66670 $D=0
M3020 325 925 921 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=52780 $D=0
M3021 326 926 922 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=57410 $D=0
M3022 327 927 923 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=62040 $D=0
M3023 328 928 924 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=66670 $D=0
M3024 925 122 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=52780 $D=0
M3025 926 122 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=57410 $D=0
M3026 927 122 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=62040 $D=0
M3027 928 122 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=66670 $D=0
M3028 191 123 929 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=52780 $D=0
M3029 192 123 930 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=57410 $D=0
M3030 193 123 931 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=62040 $D=0
M3031 194 123 932 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=66670 $D=0
M3032 933 124 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=52780 $D=0
M3033 934 124 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=57410 $D=0
M3034 935 124 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=62040 $D=0
M3035 936 124 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=66670 $D=0
M3036 8 933 317 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=52780 $D=0
M3037 9 934 318 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=57410 $D=0
M3038 10 935 319 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=62040 $D=0
M3039 11 936 320 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=66670 $D=0
M3040 325 929 8 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=52780 $D=0
M3041 326 930 9 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=57410 $D=0
M3042 327 931 10 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=62040 $D=0
M3043 328 932 11 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=66670 $D=0
M3044 191 941 937 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=52780 $D=0
M3045 192 942 938 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=57410 $D=0
M3046 193 943 939 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=62040 $D=0
M3047 194 944 940 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=66670 $D=0
M3048 941 126 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=52780 $D=0
M3049 942 126 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=57410 $D=0
M3050 943 126 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=62040 $D=0
M3051 944 126 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=66670 $D=0
M3052 1373 317 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=52780 $D=0
M3053 1374 318 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=57410 $D=0
M3054 1375 319 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=62040 $D=0
M3055 1376 320 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=66670 $D=0
M3056 945 941 1373 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=52780 $D=0
M3057 946 942 1374 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=57410 $D=0
M3058 947 943 1375 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=62040 $D=0
M3059 948 944 1376 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=66670 $D=0
M3060 191 945 949 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=52780 $D=0
M3061 192 946 950 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=57410 $D=0
M3062 193 947 951 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=62040 $D=0
M3063 194 948 952 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=66670 $D=0
M3064 1377 949 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=52780 $D=0
M3065 1378 950 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=57410 $D=0
M3066 1379 951 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=62040 $D=0
M3067 1380 952 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=66670 $D=0
M3068 945 937 1377 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=52780 $D=0
M3069 946 938 1378 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=57410 $D=0
M3070 947 939 1379 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=62040 $D=0
M3071 948 940 1380 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=66670 $D=0
M3072 191 957 953 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=52780 $D=0
M3073 192 958 954 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=57410 $D=0
M3074 193 959 955 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=62040 $D=0
M3075 194 960 956 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=66670 $D=0
M3076 957 126 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=52780 $D=0
M3077 958 126 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=57410 $D=0
M3078 959 126 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=62040 $D=0
M3079 960 126 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=66670 $D=0
M3080 1381 325 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=52780 $D=0
M3081 1382 326 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=57410 $D=0
M3082 1383 327 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=62040 $D=0
M3083 1384 328 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=66670 $D=0
M3084 961 957 1381 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=52780 $D=0
M3085 962 958 1382 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=57410 $D=0
M3086 963 959 1383 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=62040 $D=0
M3087 964 960 1384 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=66670 $D=0
M3088 191 961 127 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=52780 $D=0
M3089 192 962 128 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=57410 $D=0
M3090 193 963 129 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=62040 $D=0
M3091 194 964 130 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=66670 $D=0
M3092 1385 127 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=52780 $D=0
M3093 1386 128 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=57410 $D=0
M3094 1387 129 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=62040 $D=0
M3095 1388 130 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=66670 $D=0
M3096 961 953 1385 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=52780 $D=0
M3097 962 954 1386 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=57410 $D=0
M3098 963 955 1387 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=62040 $D=0
M3099 964 956 1388 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=66670 $D=0
M3100 965 131 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=52780 $D=0
M3101 966 131 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=57410 $D=0
M3102 967 131 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=62040 $D=0
M3103 968 131 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=66670 $D=0
M3104 969 131 949 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=52780 $D=0
M3105 970 131 950 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=57410 $D=0
M3106 971 131 951 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=62040 $D=0
M3107 972 131 952 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=66670 $D=0
M3108 132 965 969 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=52780 $D=0
M3109 132 966 970 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=57410 $D=0
M3110 132 967 971 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=62040 $D=0
M3111 132 968 972 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=66670 $D=0
M3112 973 133 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=52780 $D=0
M3113 974 133 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=57410 $D=0
M3114 975 133 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=62040 $D=0
M3115 976 133 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=66670 $D=0
M3116 977 133 127 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=52780 $D=0
M3117 978 133 128 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=57410 $D=0
M3118 979 133 129 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=62040 $D=0
M3119 980 133 130 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=66670 $D=0
M3120 1389 973 977 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=52780 $D=0
M3121 1390 974 978 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=57410 $D=0
M3122 1391 975 979 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=62040 $D=0
M3123 1392 976 980 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=66670 $D=0
M3124 191 127 1389 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=52780 $D=0
M3125 192 128 1390 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=57410 $D=0
M3126 193 129 1391 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=62040 $D=0
M3127 194 130 1392 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=66670 $D=0
M3128 981 134 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=52780 $D=0
M3129 982 134 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=57410 $D=0
M3130 983 134 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=62040 $D=0
M3131 984 134 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=66670 $D=0
M3132 985 134 977 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=52780 $D=0
M3133 986 134 978 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=57410 $D=0
M3134 987 134 979 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=62040 $D=0
M3135 988 134 980 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=66670 $D=0
M3136 15 981 985 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=52780 $D=0
M3137 16 982 986 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=57410 $D=0
M3138 17 983 987 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=62040 $D=0
M3139 18 984 988 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=66670 $D=0
M3140 992 989 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=52780 $D=0
M3141 993 990 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=57410 $D=0
M3142 994 991 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=62040 $D=0
M3143 995 135 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=66670 $D=0
M3144 191 1000 996 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=52780 $D=0
M3145 192 1001 997 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=57410 $D=0
M3146 193 1002 998 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=62040 $D=0
M3147 194 1003 999 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=66670 $D=0
M3148 1004 969 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=52780 $D=0
M3149 1005 970 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=57410 $D=0
M3150 1006 971 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=62040 $D=0
M3151 1007 972 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=66670 $D=0
M3152 1000 969 989 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=52780 $D=0
M3153 1001 970 990 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=57410 $D=0
M3154 1002 971 991 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=62040 $D=0
M3155 1003 972 135 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=66670 $D=0
M3156 992 1004 1000 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=52780 $D=0
M3157 993 1005 1001 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=57410 $D=0
M3158 994 1006 1002 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=62040 $D=0
M3159 995 1007 1003 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=66670 $D=0
M3160 1008 996 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=52780 $D=0
M3161 1009 997 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=57410 $D=0
M3162 1010 998 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=62040 $D=0
M3163 1011 999 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=66670 $D=0
M3164 136 996 985 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=52780 $D=0
M3165 989 997 986 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=57410 $D=0
M3166 990 998 987 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=62040 $D=0
M3167 991 999 988 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=66670 $D=0
M3168 969 1008 136 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=52780 $D=0
M3169 970 1009 989 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=57410 $D=0
M3170 971 1010 990 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=62040 $D=0
M3171 972 1011 991 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=66670 $D=0
M3172 1012 136 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=52780 $D=0
M3173 1013 989 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=57410 $D=0
M3174 1014 990 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=62040 $D=0
M3175 1015 991 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=66670 $D=0
M3176 1016 996 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=52780 $D=0
M3177 1017 997 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=57410 $D=0
M3178 1018 998 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=62040 $D=0
M3179 1019 999 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=66670 $D=0
M3180 1020 996 1012 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=52780 $D=0
M3181 1021 997 1013 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=57410 $D=0
M3182 1022 998 1014 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=62040 $D=0
M3183 1023 999 1015 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=66670 $D=0
M3184 985 1016 1020 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=52780 $D=0
M3185 986 1017 1021 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=57410 $D=0
M3186 987 1018 1022 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=62040 $D=0
M3187 988 1019 1023 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=66670 $D=0
M3188 1413 969 191 191 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=52420 $D=0
M3189 1414 970 192 192 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=57050 $D=0
M3190 1415 971 193 193 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=61680 $D=0
M3191 1416 972 194 194 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=66310 $D=0
M3192 1024 985 1413 191 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=52420 $D=0
M3193 1025 986 1414 192 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=57050 $D=0
M3194 1026 987 1415 193 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=61680 $D=0
M3195 1027 988 1416 194 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=66310 $D=0
M3196 1028 1020 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=52780 $D=0
M3197 1029 1021 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=57410 $D=0
M3198 1030 1022 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=62040 $D=0
M3199 1031 1023 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=66670 $D=0
M3200 1032 969 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=52780 $D=0
M3201 1033 970 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=57410 $D=0
M3202 1034 971 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=62040 $D=0
M3203 1035 972 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=66670 $D=0
M3204 191 985 1032 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=52780 $D=0
M3205 192 986 1033 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=57410 $D=0
M3206 193 987 1034 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=62040 $D=0
M3207 194 988 1035 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=66670 $D=0
M3208 1036 969 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=52780 $D=0
M3209 1037 970 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=57410 $D=0
M3210 1038 971 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=62040 $D=0
M3211 1039 972 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=66670 $D=0
M3212 191 985 1036 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=52780 $D=0
M3213 192 986 1037 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=57410 $D=0
M3214 193 987 1038 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=62040 $D=0
M3215 194 988 1039 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=66670 $D=0
M3216 1417 969 191 191 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=52600 $D=0
M3217 1418 970 192 192 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=57230 $D=0
M3218 1419 971 193 193 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=61860 $D=0
M3219 1420 972 194 194 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=66490 $D=0
M3220 1044 985 1417 191 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=52600 $D=0
M3221 1045 986 1418 192 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=57230 $D=0
M3222 1046 987 1419 193 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=61860 $D=0
M3223 1047 988 1420 194 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=66490 $D=0
M3224 191 1036 1044 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=52780 $D=0
M3225 192 1037 1045 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=57410 $D=0
M3226 193 1038 1046 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=62040 $D=0
M3227 194 1039 1047 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=66670 $D=0
M3228 1048 140 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=52780 $D=0
M3229 1049 140 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=57410 $D=0
M3230 1050 140 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=62040 $D=0
M3231 1051 140 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=66670 $D=0
M3232 1052 140 1024 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=52780 $D=0
M3233 1053 140 1025 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=57410 $D=0
M3234 1054 140 1026 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=62040 $D=0
M3235 1055 140 1027 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=66670 $D=0
M3236 1032 1048 1052 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=52780 $D=0
M3237 1033 1049 1053 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=57410 $D=0
M3238 1034 1050 1054 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=62040 $D=0
M3239 1035 1051 1055 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=66670 $D=0
M3240 1056 140 1028 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=52780 $D=0
M3241 1057 140 1029 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=57410 $D=0
M3242 1058 140 1030 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=62040 $D=0
M3243 1059 140 1031 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=66670 $D=0
M3244 1044 1048 1056 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=52780 $D=0
M3245 1045 1049 1057 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=57410 $D=0
M3246 1046 1050 1058 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=62040 $D=0
M3247 1047 1051 1059 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=66670 $D=0
M3248 1060 141 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=52780 $D=0
M3249 1061 141 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=57410 $D=0
M3250 1062 141 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=62040 $D=0
M3251 1063 141 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=66670 $D=0
M3252 1064 141 1056 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=52780 $D=0
M3253 1065 141 1057 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=57410 $D=0
M3254 1066 141 1058 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=62040 $D=0
M3255 1067 141 1059 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=66670 $D=0
M3256 1052 1060 1064 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=52780 $D=0
M3257 1053 1061 1065 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=57410 $D=0
M3258 1054 1062 1066 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=62040 $D=0
M3259 1055 1063 1067 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=66670 $D=0
M3260 19 1064 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=52780 $D=0
M3261 20 1065 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=57410 $D=0
M3262 21 1066 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=62040 $D=0
M3263 22 1067 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=66670 $D=0
M3264 1068 142 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=52780 $D=0
M3265 1069 142 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=57410 $D=0
M3266 1070 142 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=62040 $D=0
M3267 1071 142 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=66670 $D=0
M3268 1072 142 143 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=52780 $D=0
M3269 1073 142 144 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=57410 $D=0
M3270 1074 142 145 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=62040 $D=0
M3271 1075 142 146 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=66670 $D=0
M3272 147 1068 1072 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=52780 $D=0
M3273 148 1069 1073 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=57410 $D=0
M3274 143 1070 1074 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=62040 $D=0
M3275 144 1071 1075 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=66670 $D=0
M3276 1076 142 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=52780 $D=0
M3277 1077 142 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=57410 $D=0
M3278 1078 142 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=62040 $D=0
M3279 1079 142 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=66670 $D=0
M3280 1080 142 149 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=52780 $D=0
M3281 1081 142 150 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=57410 $D=0
M3282 1082 142 151 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=62040 $D=0
M3283 1083 142 152 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=66670 $D=0
M3284 153 1076 1080 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=52780 $D=0
M3285 154 1077 1081 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=57410 $D=0
M3286 155 1078 1082 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=62040 $D=0
M3287 156 1079 1083 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=66670 $D=0
M3288 1084 142 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=52780 $D=0
M3289 1085 142 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=57410 $D=0
M3290 1086 142 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=62040 $D=0
M3291 1087 142 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=66670 $D=0
M3292 1088 142 137 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=52780 $D=0
M3293 1089 142 139 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=57410 $D=0
M3294 1090 142 138 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=62040 $D=0
M3295 1091 142 157 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=66670 $D=0
M3296 158 1084 1088 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=52780 $D=0
M3297 120 1085 1089 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=57410 $D=0
M3298 121 1086 1090 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=62040 $D=0
M3299 125 1087 1091 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=66670 $D=0
M3300 1092 142 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=52780 $D=0
M3301 1093 142 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=57410 $D=0
M3302 1094 142 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=62040 $D=0
M3303 1095 142 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=66670 $D=0
M3304 1096 142 159 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=52780 $D=0
M3305 1097 142 160 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=57410 $D=0
M3306 1098 142 161 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=62040 $D=0
M3307 1099 142 162 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=66670 $D=0
M3308 163 1092 1096 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=52780 $D=0
M3309 164 1093 1097 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=57410 $D=0
M3310 165 1094 1098 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=62040 $D=0
M3311 166 1095 1099 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=66670 $D=0
M3312 1100 142 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=52780 $D=0
M3313 1101 142 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=57410 $D=0
M3314 1102 142 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=62040 $D=0
M3315 1103 142 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=66670 $D=0
M3316 1104 142 167 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=52780 $D=0
M3317 1105 142 168 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=57410 $D=0
M3318 1106 142 169 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=62040 $D=0
M3319 1107 142 170 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=66670 $D=0
M3320 171 1100 1104 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=52780 $D=0
M3321 171 1101 1105 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=57410 $D=0
M3322 171 1102 1106 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=62040 $D=0
M3323 171 1103 1107 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=66670 $D=0
M3324 191 969 1393 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=52780 $D=0
M3325 192 970 1394 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=57410 $D=0
M3326 193 971 1395 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=62040 $D=0
M3327 194 972 1396 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=66670 $D=0
M3328 148 1393 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=52780 $D=0
M3329 143 1394 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=57410 $D=0
M3330 144 1395 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=62040 $D=0
M3331 145 1396 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=66670 $D=0
M3332 1108 172 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=52780 $D=0
M3333 1109 172 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=57410 $D=0
M3334 1110 172 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=62040 $D=0
M3335 1111 172 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=66670 $D=0
M3336 155 172 148 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=52780 $D=0
M3337 156 172 143 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=57410 $D=0
M3338 149 172 144 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=62040 $D=0
M3339 150 172 145 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=66670 $D=0
M3340 1072 1108 155 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=52780 $D=0
M3341 1073 1109 156 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=57410 $D=0
M3342 1074 1110 149 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=62040 $D=0
M3343 1075 1111 150 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=66670 $D=0
M3344 1112 173 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=52780 $D=0
M3345 1113 173 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=57410 $D=0
M3346 1114 173 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=62040 $D=0
M3347 1115 173 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=66670 $D=0
M3348 174 173 155 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=52780 $D=0
M3349 114 173 156 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=57410 $D=0
M3350 115 173 149 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=62040 $D=0
M3351 119 173 150 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=66670 $D=0
M3352 1080 1112 174 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=52780 $D=0
M3353 1081 1113 114 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=57410 $D=0
M3354 1082 1114 115 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=62040 $D=0
M3355 1083 1115 119 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=66670 $D=0
M3356 1116 175 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=52780 $D=0
M3357 1117 175 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=57410 $D=0
M3358 1118 175 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=62040 $D=0
M3359 1119 175 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=66670 $D=0
M3360 174 175 174 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=52780 $D=0
M3361 114 175 114 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=57410 $D=0
M3362 115 175 115 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=62040 $D=0
M3363 119 175 119 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=66670 $D=0
M3364 1088 1116 174 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=52780 $D=0
M3365 1089 1117 114 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=57410 $D=0
M3366 1090 1118 115 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=62040 $D=0
M3367 1091 1119 119 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=66670 $D=0
M3368 1120 176 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=52780 $D=0
M3369 1121 176 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=57410 $D=0
M3370 1122 176 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=62040 $D=0
M3371 1123 176 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=66670 $D=0
M3372 177 176 174 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=52780 $D=0
M3373 178 176 114 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=57410 $D=0
M3374 179 176 115 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=62040 $D=0
M3375 180 176 119 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=66670 $D=0
M3376 1096 1120 177 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=52780 $D=0
M3377 1097 1121 178 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=57410 $D=0
M3378 1098 1122 179 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=62040 $D=0
M3379 1099 1123 180 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=66670 $D=0
M3380 1124 181 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=52780 $D=0
M3381 1125 181 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=57410 $D=0
M3382 1126 181 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=62040 $D=0
M3383 1127 181 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=66670 $D=0
M3384 269 181 177 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=52780 $D=0
M3385 270 181 178 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=57410 $D=0
M3386 271 181 179 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=62040 $D=0
M3387 272 181 180 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=66670 $D=0
M3388 1104 1124 269 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=52780 $D=0
M3389 1105 1125 270 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=57410 $D=0
M3390 1106 1126 271 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=62040 $D=0
M3391 1107 1127 272 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=66670 $D=0
M3392 1128 182 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=52780 $D=0
M3393 1129 182 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=57410 $D=0
M3394 1130 182 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=62040 $D=0
M3395 1131 182 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=66670 $D=0
M3396 1132 182 127 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=52780 $D=0
M3397 1133 182 128 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=57410 $D=0
M3398 1134 182 129 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=62040 $D=0
M3399 1135 182 130 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=66670 $D=0
M3400 15 1128 1132 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=52780 $D=0
M3401 16 1129 1133 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=57410 $D=0
M3402 17 1130 1134 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=62040 $D=0
M3403 18 1131 1135 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=66670 $D=0
M3404 1136 949 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=52780 $D=0
M3405 1137 950 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=57410 $D=0
M3406 1138 951 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=62040 $D=0
M3407 1139 952 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=66670 $D=0
M3408 191 1132 1136 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=52780 $D=0
M3409 192 1133 1137 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=57410 $D=0
M3410 193 1134 1138 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=62040 $D=0
M3411 194 1135 1139 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=66670 $D=0
M3412 1421 949 191 191 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=52600 $D=0
M3413 1422 950 192 192 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=57230 $D=0
M3414 1423 951 193 193 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=61860 $D=0
M3415 1424 952 194 194 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=66490 $D=0
M3416 1144 1132 1421 191 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=52600 $D=0
M3417 1145 1133 1422 192 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=57230 $D=0
M3418 1146 1134 1423 193 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=61860 $D=0
M3419 1147 1135 1424 194 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=66490 $D=0
M3420 191 1136 1144 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=52780 $D=0
M3421 192 1137 1145 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=57410 $D=0
M3422 193 1138 1146 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=62040 $D=0
M3423 194 1139 1147 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=66670 $D=0
M3424 1397 183 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=52780 $D=0
M3425 1398 1148 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=57410 $D=0
M3426 1399 1149 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=62040 $D=0
M3427 1400 1150 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=66670 $D=0
M3428 191 1144 1397 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=52780 $D=0
M3429 192 1145 1398 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=57410 $D=0
M3430 193 1146 1399 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=62040 $D=0
M3431 194 1147 1400 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=66670 $D=0
M3432 1148 1397 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=52780 $D=0
M3433 1149 1398 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=57410 $D=0
M3434 1150 1399 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=62040 $D=0
M3435 184 1400 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=66670 $D=0
M3436 1425 949 191 191 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=52420 $D=0
M3437 1426 950 192 192 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=57050 $D=0
M3438 1427 951 193 193 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=61680 $D=0
M3439 1428 952 194 194 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=66310 $D=0
M3440 1151 1155 1425 191 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=52420 $D=0
M3441 1152 1156 1426 192 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=57050 $D=0
M3442 1153 1157 1427 193 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=61680 $D=0
M3443 1154 1158 1428 194 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=66310 $D=0
M3444 1155 1132 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=52780 $D=0
M3445 1156 1133 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=57410 $D=0
M3446 1157 1134 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=62040 $D=0
M3447 1158 1135 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=66670 $D=0
M3448 1159 1151 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=52780 $D=0
M3449 1160 1152 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=57410 $D=0
M3450 1161 1153 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=62040 $D=0
M3451 1162 1154 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=66670 $D=0
M3452 191 183 1159 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=52780 $D=0
M3453 192 1148 1160 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=57410 $D=0
M3454 193 1149 1161 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=62040 $D=0
M3455 194 1150 1162 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=66670 $D=0
M3456 1166 185 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=52780 $D=0
M3457 1167 1163 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=57410 $D=0
M3458 1168 1164 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=62040 $D=0
M3459 1169 1165 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=66670 $D=0
M3460 1163 1159 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=52780 $D=0
M3461 1164 1160 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=57410 $D=0
M3462 1165 1161 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=62040 $D=0
M3463 186 1162 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=66670 $D=0
M3464 191 1166 1163 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=52780 $D=0
M3465 192 1167 1164 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=57410 $D=0
M3466 193 1168 1165 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=62040 $D=0
M3467 194 1169 186 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=66670 $D=0
M3468 1173 1170 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=52780 $D=0
M3469 1174 1171 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=57410 $D=0
M3470 1175 1172 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=62040 $D=0
M3471 1176 187 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=66670 $D=0
M3472 191 1181 1177 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=52780 $D=0
M3473 192 1182 1178 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=57410 $D=0
M3474 193 1183 1179 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=62040 $D=0
M3475 194 1184 1180 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=66670 $D=0
M3476 1185 132 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=52780 $D=0
M3477 1186 132 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=57410 $D=0
M3478 1187 132 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=62040 $D=0
M3479 1188 132 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=66670 $D=0
M3480 1181 132 1170 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=52780 $D=0
M3481 1182 132 1171 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=57410 $D=0
M3482 1183 132 1172 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=62040 $D=0
M3483 1184 132 187 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=66670 $D=0
M3484 1173 1185 1181 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=52780 $D=0
M3485 1174 1186 1182 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=57410 $D=0
M3486 1175 1187 1183 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=62040 $D=0
M3487 1176 1188 1184 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=66670 $D=0
M3488 1189 1177 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=52780 $D=0
M3489 1190 1178 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=57410 $D=0
M3490 1191 1179 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=62040 $D=0
M3491 1192 1180 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=66670 $D=0
M3492 188 1177 8 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=52780 $D=0
M3493 1170 1178 9 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=57410 $D=0
M3494 1171 1179 10 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=62040 $D=0
M3495 1172 1180 11 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=66670 $D=0
M3496 132 1189 188 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=52780 $D=0
M3497 132 1190 1170 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=57410 $D=0
M3498 132 1191 1171 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=62040 $D=0
M3499 132 1192 1172 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=66670 $D=0
M3500 1193 188 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=52780 $D=0
M3501 1194 1170 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=57410 $D=0
M3502 1195 1171 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=62040 $D=0
M3503 1196 1172 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=66670 $D=0
M3504 1197 1177 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=52780 $D=0
M3505 1198 1178 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=57410 $D=0
M3506 1199 1179 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=62040 $D=0
M3507 1200 1180 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=66670 $D=0
M3508 273 1177 1193 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=52780 $D=0
M3509 274 1178 1194 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=57410 $D=0
M3510 275 1179 1195 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=62040 $D=0
M3511 276 1180 1196 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=66670 $D=0
M3512 8 1197 273 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=52780 $D=0
M3513 9 1198 274 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=57410 $D=0
M3514 10 1199 275 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=62040 $D=0
M3515 11 1200 276 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=66670 $D=0
M3516 1201 189 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=52780 $D=0
M3517 1202 189 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=57410 $D=0
M3518 1203 189 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=62040 $D=0
M3519 1204 189 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=66670 $D=0
M3520 1205 189 273 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=52780 $D=0
M3521 1206 189 274 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=57410 $D=0
M3522 1207 189 275 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=62040 $D=0
M3523 1208 189 276 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=66670 $D=0
M3524 19 1201 1205 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=52780 $D=0
M3525 20 1202 1206 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=57410 $D=0
M3526 21 1203 1207 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=62040 $D=0
M3527 22 1204 1208 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=66670 $D=0
M3528 1209 190 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=52780 $D=0
M3529 1210 190 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=57410 $D=0
M3530 1211 190 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=62040 $D=0
M3531 1212 190 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=66670 $D=0
M3532 190 190 1205 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=52780 $D=0
M3533 190 190 1206 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=57410 $D=0
M3534 190 190 1207 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=62040 $D=0
M3535 190 190 1208 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=66670 $D=0
M3536 8 1209 190 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=52780 $D=0
M3537 9 1210 190 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=57410 $D=0
M3538 10 1211 190 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=62040 $D=0
M3539 11 1212 190 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=66670 $D=0
M3540 1213 126 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=52780 $D=0
M3541 1214 126 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=57410 $D=0
M3542 1215 126 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=62040 $D=0
M3543 1216 126 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=66670 $D=0
M3544 191 1213 1217 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=52780 $D=0
M3545 192 1214 1218 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=57410 $D=0
M3546 193 1215 1219 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=62040 $D=0
M3547 194 1216 1220 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=66670 $D=0
M3548 1221 126 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=52780 $D=0
M3549 1222 126 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=57410 $D=0
M3550 1223 126 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=62040 $D=0
M3551 1224 126 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=66670 $D=0
M3552 1225 1217 190 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=52780 $D=0
M3553 1226 1218 190 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=57410 $D=0
M3554 1227 1219 190 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=62040 $D=0
M3555 1228 1220 190 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=66670 $D=0
M3556 191 1225 1401 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=52780 $D=0
M3557 192 1226 1402 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=57410 $D=0
M3558 193 1227 1403 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=62040 $D=0
M3559 194 1228 1404 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=66670 $D=0
M3560 1229 1401 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=52780 $D=0
M3561 1230 1402 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=57410 $D=0
M3562 1231 1403 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=62040 $D=0
M3563 1232 1404 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=66670 $D=0
M3564 1225 1213 1229 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=52780 $D=0
M3565 1226 1214 1230 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=57410 $D=0
M3566 1227 1215 1231 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=62040 $D=0
M3567 1228 1216 1232 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=66670 $D=0
M3568 1233 1221 1229 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=52780 $D=0
M3569 1234 1222 1230 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=57410 $D=0
M3570 1235 1223 1231 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=62040 $D=0
M3571 1236 1224 1232 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=66670 $D=0
M3572 191 1241 1237 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=52780 $D=0
M3573 192 1242 1238 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=57410 $D=0
M3574 193 1243 1239 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=62040 $D=0
M3575 194 1244 1240 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=66670 $D=0
M3576 1241 126 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=52780 $D=0
M3577 1242 126 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=57410 $D=0
M3578 1243 126 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=62040 $D=0
M3579 1244 126 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=66670 $D=0
M3580 1405 1233 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=52780 $D=0
M3581 1406 1234 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=57410 $D=0
M3582 1407 1235 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=62040 $D=0
M3583 1408 1236 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=66670 $D=0
M3584 1245 1241 1405 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=52780 $D=0
M3585 1246 1242 1406 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=57410 $D=0
M3586 1247 1243 1407 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=62040 $D=0
M3587 1248 1244 1408 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=66670 $D=0
M3588 191 1245 132 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=52780 $D=0
M3589 192 1246 132 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=57410 $D=0
M3590 193 1247 132 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=62040 $D=0
M3591 194 1248 132 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=66670 $D=0
M3592 1409 132 191 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=52780 $D=0
M3593 1410 132 192 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=57410 $D=0
M3594 1411 132 193 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=62040 $D=0
M3595 1412 132 194 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=66670 $D=0
M3596 1245 1237 1409 191 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=52780 $D=0
M3597 1246 1238 1410 192 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=57410 $D=0
M3598 1247 1239 1411 193 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=62040 $D=0
M3599 1248 1240 1412 194 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=66670 $D=0
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 109 110 111 112 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166
** N=811 EP=163 IP=1514 FDC=1800
M0 197 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=42270 $D=1
M1 198 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=46900 $D=1
M2 199 197 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=42270 $D=1
M3 200 198 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=46900 $D=1
M4 6 1 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=42270 $D=1
M5 7 1 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=46900 $D=1
M6 201 197 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=42270 $D=1
M7 202 198 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=46900 $D=1
M8 5 1 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=42270 $D=1
M9 5 1 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=46900 $D=1
M10 203 197 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=42270 $D=1
M11 204 198 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=46900 $D=1
M12 6 1 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=42270 $D=1
M13 7 1 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=46900 $D=1
M14 207 205 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=42270 $D=1
M15 208 206 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=46900 $D=1
M16 205 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=42270 $D=1
M17 206 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=46900 $D=1
M18 209 205 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=42270 $D=1
M19 210 206 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=46900 $D=1
M20 199 9 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=42270 $D=1
M21 200 9 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=46900 $D=1
M22 211 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=42270 $D=1
M23 212 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=46900 $D=1
M24 213 211 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=42270 $D=1
M25 214 212 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=46900 $D=1
M26 207 10 213 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=42270 $D=1
M27 208 10 214 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=46900 $D=1
M28 215 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=42270 $D=1
M29 216 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=46900 $D=1
M30 217 215 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=42270 $D=1
M31 218 216 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=46900 $D=1
M32 12 11 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=42270 $D=1
M33 13 11 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=46900 $D=1
M34 219 215 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=42270 $D=1
M35 220 216 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=46900 $D=1
M36 221 11 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=42270 $D=1
M37 222 11 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=46900 $D=1
M38 225 215 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=42270 $D=1
M39 226 216 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=46900 $D=1
M40 213 11 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=42270 $D=1
M41 214 11 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=46900 $D=1
M42 229 227 225 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=42270 $D=1
M43 230 228 226 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=46900 $D=1
M44 227 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=42270 $D=1
M45 228 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=46900 $D=1
M46 231 227 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=42270 $D=1
M47 232 228 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=46900 $D=1
M48 217 16 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=42270 $D=1
M49 218 16 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=46900 $D=1
M50 233 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=42270 $D=1
M51 234 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=46900 $D=1
M52 235 233 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=42270 $D=1
M53 236 234 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=46900 $D=1
M54 229 17 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=42270 $D=1
M55 230 17 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=46900 $D=1
M56 6 18 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=42270 $D=1
M57 7 18 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=46900 $D=1
M58 239 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=42270 $D=1
M59 240 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=46900 $D=1
M60 241 18 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=42270 $D=1
M61 242 18 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=46900 $D=1
M62 6 241 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=42270 $D=1
M63 7 242 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=46900 $D=1
M64 243 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=42270 $D=1
M65 244 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=46900 $D=1
M66 241 237 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=42270 $D=1
M67 242 238 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=46900 $D=1
M68 243 19 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=42270 $D=1
M69 244 19 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=46900 $D=1
M70 249 20 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=42270 $D=1
M71 250 20 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=46900 $D=1
M72 247 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=42270 $D=1
M73 248 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=46900 $D=1
M74 6 21 251 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=42270 $D=1
M75 7 21 252 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=46900 $D=1
M76 253 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=42270 $D=1
M77 254 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=46900 $D=1
M78 255 21 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=42270 $D=1
M79 256 21 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=46900 $D=1
M80 6 255 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=42270 $D=1
M81 7 256 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=46900 $D=1
M82 257 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=42270 $D=1
M83 258 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=46900 $D=1
M84 255 251 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=42270 $D=1
M85 256 252 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=46900 $D=1
M86 257 22 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=42270 $D=1
M87 258 22 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=46900 $D=1
M88 249 23 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=42270 $D=1
M89 250 23 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=46900 $D=1
M90 259 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=42270 $D=1
M91 260 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=46900 $D=1
M92 6 24 261 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=42270 $D=1
M93 7 24 262 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=46900 $D=1
M94 263 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=42270 $D=1
M95 264 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=46900 $D=1
M96 265 24 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=42270 $D=1
M97 266 24 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=46900 $D=1
M98 6 265 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=42270 $D=1
M99 7 266 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=46900 $D=1
M100 267 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=42270 $D=1
M101 268 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=46900 $D=1
M102 265 261 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=42270 $D=1
M103 266 262 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=46900 $D=1
M104 267 25 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=42270 $D=1
M105 268 25 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=46900 $D=1
M106 249 26 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=42270 $D=1
M107 250 26 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=46900 $D=1
M108 269 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=42270 $D=1
M109 270 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=46900 $D=1
M110 6 27 271 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=42270 $D=1
M111 7 27 272 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=46900 $D=1
M112 273 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=42270 $D=1
M113 274 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=46900 $D=1
M114 275 27 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=42270 $D=1
M115 276 27 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=46900 $D=1
M116 6 275 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=42270 $D=1
M117 7 276 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=46900 $D=1
M118 277 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=42270 $D=1
M119 278 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=46900 $D=1
M120 275 271 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=42270 $D=1
M121 276 272 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=46900 $D=1
M122 277 28 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=42270 $D=1
M123 278 28 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=46900 $D=1
M124 249 29 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=42270 $D=1
M125 250 29 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=46900 $D=1
M126 279 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=42270 $D=1
M127 280 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=46900 $D=1
M128 6 30 281 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=42270 $D=1
M129 7 30 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=46900 $D=1
M130 283 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=42270 $D=1
M131 284 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=46900 $D=1
M132 285 30 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=42270 $D=1
M133 286 30 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=46900 $D=1
M134 6 285 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=42270 $D=1
M135 7 286 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=46900 $D=1
M136 287 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=42270 $D=1
M137 288 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=46900 $D=1
M138 285 281 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=42270 $D=1
M139 286 282 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=46900 $D=1
M140 287 31 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=42270 $D=1
M141 288 31 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=46900 $D=1
M142 249 32 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=42270 $D=1
M143 250 32 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=46900 $D=1
M144 289 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=42270 $D=1
M145 290 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=46900 $D=1
M146 6 33 291 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=42270 $D=1
M147 7 33 292 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=46900 $D=1
M148 293 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=42270 $D=1
M149 294 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=46900 $D=1
M150 295 33 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=42270 $D=1
M151 296 33 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=46900 $D=1
M152 6 295 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=42270 $D=1
M153 7 296 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=46900 $D=1
M154 297 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=42270 $D=1
M155 298 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=46900 $D=1
M156 295 291 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=42270 $D=1
M157 296 292 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=46900 $D=1
M158 297 34 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=42270 $D=1
M159 298 34 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=46900 $D=1
M160 249 35 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=42270 $D=1
M161 250 35 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=46900 $D=1
M162 299 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=42270 $D=1
M163 300 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=46900 $D=1
M164 6 36 301 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=42270 $D=1
M165 7 36 302 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=46900 $D=1
M166 303 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=42270 $D=1
M167 304 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=46900 $D=1
M168 305 36 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=42270 $D=1
M169 306 36 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=46900 $D=1
M170 6 305 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=42270 $D=1
M171 7 306 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=46900 $D=1
M172 307 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=42270 $D=1
M173 308 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=46900 $D=1
M174 305 301 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=42270 $D=1
M175 306 302 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=46900 $D=1
M176 307 37 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=42270 $D=1
M177 308 37 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=46900 $D=1
M178 249 38 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=42270 $D=1
M179 250 38 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=46900 $D=1
M180 309 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=42270 $D=1
M181 310 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=46900 $D=1
M182 6 39 311 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=42270 $D=1
M183 7 39 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=46900 $D=1
M184 313 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=42270 $D=1
M185 314 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=46900 $D=1
M186 315 39 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=42270 $D=1
M187 316 39 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=46900 $D=1
M188 6 315 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=42270 $D=1
M189 7 316 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=46900 $D=1
M190 317 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=42270 $D=1
M191 318 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=46900 $D=1
M192 315 311 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=42270 $D=1
M193 316 312 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=46900 $D=1
M194 317 40 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=42270 $D=1
M195 318 40 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=46900 $D=1
M196 249 41 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=42270 $D=1
M197 250 41 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=46900 $D=1
M198 319 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=42270 $D=1
M199 320 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=46900 $D=1
M200 6 42 321 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=42270 $D=1
M201 7 42 322 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=46900 $D=1
M202 323 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=42270 $D=1
M203 324 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=46900 $D=1
M204 325 42 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=42270 $D=1
M205 326 42 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=46900 $D=1
M206 6 325 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=42270 $D=1
M207 7 326 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=46900 $D=1
M208 327 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=42270 $D=1
M209 328 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=46900 $D=1
M210 325 321 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=42270 $D=1
M211 326 322 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=46900 $D=1
M212 327 43 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=42270 $D=1
M213 328 43 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=46900 $D=1
M214 249 44 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=42270 $D=1
M215 250 44 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=46900 $D=1
M216 329 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=42270 $D=1
M217 330 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=46900 $D=1
M218 6 45 331 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=42270 $D=1
M219 7 45 332 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=46900 $D=1
M220 333 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=42270 $D=1
M221 334 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=46900 $D=1
M222 335 45 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=42270 $D=1
M223 336 45 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=46900 $D=1
M224 6 335 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=42270 $D=1
M225 7 336 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=46900 $D=1
M226 337 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=42270 $D=1
M227 338 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=46900 $D=1
M228 335 331 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=42270 $D=1
M229 336 332 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=46900 $D=1
M230 337 46 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=42270 $D=1
M231 338 46 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=46900 $D=1
M232 249 47 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=42270 $D=1
M233 250 47 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=46900 $D=1
M234 339 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=42270 $D=1
M235 340 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=46900 $D=1
M236 6 48 341 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=42270 $D=1
M237 7 48 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=46900 $D=1
M238 343 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=42270 $D=1
M239 344 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=46900 $D=1
M240 345 48 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=42270 $D=1
M241 346 48 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=46900 $D=1
M242 6 345 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=42270 $D=1
M243 7 346 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=46900 $D=1
M244 347 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=42270 $D=1
M245 348 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=46900 $D=1
M246 345 341 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=42270 $D=1
M247 346 342 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=46900 $D=1
M248 347 49 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=42270 $D=1
M249 348 49 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=46900 $D=1
M250 249 50 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=42270 $D=1
M251 250 50 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=46900 $D=1
M252 349 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=42270 $D=1
M253 350 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=46900 $D=1
M254 6 51 351 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=42270 $D=1
M255 7 51 352 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=46900 $D=1
M256 353 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=42270 $D=1
M257 354 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=46900 $D=1
M258 355 51 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=42270 $D=1
M259 356 51 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=46900 $D=1
M260 6 355 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=42270 $D=1
M261 7 356 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=46900 $D=1
M262 357 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=42270 $D=1
M263 358 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=46900 $D=1
M264 355 351 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=42270 $D=1
M265 356 352 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=46900 $D=1
M266 357 52 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=42270 $D=1
M267 358 52 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=46900 $D=1
M268 249 53 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=42270 $D=1
M269 250 53 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=46900 $D=1
M270 359 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=42270 $D=1
M271 360 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=46900 $D=1
M272 6 54 361 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=42270 $D=1
M273 7 54 362 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=46900 $D=1
M274 363 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=42270 $D=1
M275 364 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=46900 $D=1
M276 365 54 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=42270 $D=1
M277 366 54 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=46900 $D=1
M278 6 365 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=42270 $D=1
M279 7 366 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=46900 $D=1
M280 367 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=42270 $D=1
M281 368 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=46900 $D=1
M282 365 361 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=42270 $D=1
M283 366 362 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=46900 $D=1
M284 367 55 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=42270 $D=1
M285 368 55 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=46900 $D=1
M286 249 56 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=42270 $D=1
M287 250 56 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=46900 $D=1
M288 369 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=42270 $D=1
M289 370 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=46900 $D=1
M290 6 57 371 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=42270 $D=1
M291 7 57 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=46900 $D=1
M292 373 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=42270 $D=1
M293 374 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=46900 $D=1
M294 375 57 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=42270 $D=1
M295 376 57 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=46900 $D=1
M296 6 375 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=42270 $D=1
M297 7 376 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=46900 $D=1
M298 377 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=42270 $D=1
M299 378 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=46900 $D=1
M300 375 371 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=42270 $D=1
M301 376 372 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=46900 $D=1
M302 377 58 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=42270 $D=1
M303 378 58 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=46900 $D=1
M304 249 59 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=42270 $D=1
M305 250 59 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=46900 $D=1
M306 379 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=42270 $D=1
M307 380 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=46900 $D=1
M308 6 60 381 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=42270 $D=1
M309 7 60 382 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=46900 $D=1
M310 383 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=42270 $D=1
M311 384 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=46900 $D=1
M312 385 60 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=42270 $D=1
M313 386 60 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=46900 $D=1
M314 6 385 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=42270 $D=1
M315 7 386 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=46900 $D=1
M316 387 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=42270 $D=1
M317 388 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=46900 $D=1
M318 385 381 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=42270 $D=1
M319 386 382 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=46900 $D=1
M320 387 61 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=42270 $D=1
M321 388 61 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=46900 $D=1
M322 249 62 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=42270 $D=1
M323 250 62 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=46900 $D=1
M324 389 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=42270 $D=1
M325 390 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=46900 $D=1
M326 6 63 391 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=42270 $D=1
M327 7 63 392 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=46900 $D=1
M328 393 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=42270 $D=1
M329 394 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=46900 $D=1
M330 395 63 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=42270 $D=1
M331 396 63 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=46900 $D=1
M332 6 395 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=42270 $D=1
M333 7 396 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=46900 $D=1
M334 397 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=42270 $D=1
M335 398 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=46900 $D=1
M336 395 391 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=42270 $D=1
M337 396 392 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=46900 $D=1
M338 397 64 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=42270 $D=1
M339 398 64 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=46900 $D=1
M340 249 65 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=42270 $D=1
M341 250 65 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=46900 $D=1
M342 399 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=42270 $D=1
M343 400 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=46900 $D=1
M344 6 66 401 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=42270 $D=1
M345 7 66 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=46900 $D=1
M346 403 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=42270 $D=1
M347 404 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=46900 $D=1
M348 405 66 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=42270 $D=1
M349 406 66 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=46900 $D=1
M350 6 405 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=42270 $D=1
M351 7 406 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=46900 $D=1
M352 407 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=42270 $D=1
M353 408 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=46900 $D=1
M354 405 401 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=42270 $D=1
M355 406 402 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=46900 $D=1
M356 407 67 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=42270 $D=1
M357 408 67 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=46900 $D=1
M358 249 68 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=42270 $D=1
M359 250 68 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=46900 $D=1
M360 409 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=42270 $D=1
M361 410 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=46900 $D=1
M362 6 69 411 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=42270 $D=1
M363 7 69 412 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=46900 $D=1
M364 413 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=42270 $D=1
M365 414 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=46900 $D=1
M366 415 69 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=42270 $D=1
M367 416 69 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=46900 $D=1
M368 6 415 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=42270 $D=1
M369 7 416 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=46900 $D=1
M370 417 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=42270 $D=1
M371 418 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=46900 $D=1
M372 415 411 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=42270 $D=1
M373 416 412 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=46900 $D=1
M374 417 70 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=42270 $D=1
M375 418 70 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=46900 $D=1
M376 249 71 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=42270 $D=1
M377 250 71 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=46900 $D=1
M378 419 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=42270 $D=1
M379 420 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=46900 $D=1
M380 6 72 421 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=42270 $D=1
M381 7 72 422 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=46900 $D=1
M382 423 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=42270 $D=1
M383 424 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=46900 $D=1
M384 425 72 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=42270 $D=1
M385 426 72 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=46900 $D=1
M386 6 425 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=42270 $D=1
M387 7 426 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=46900 $D=1
M388 427 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=42270 $D=1
M389 428 747 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=46900 $D=1
M390 425 421 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=42270 $D=1
M391 426 422 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=46900 $D=1
M392 427 73 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=42270 $D=1
M393 428 73 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=46900 $D=1
M394 249 74 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=42270 $D=1
M395 250 74 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=46900 $D=1
M396 429 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=42270 $D=1
M397 430 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=46900 $D=1
M398 6 75 431 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=42270 $D=1
M399 7 75 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=46900 $D=1
M400 433 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=42270 $D=1
M401 434 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=46900 $D=1
M402 435 75 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=42270 $D=1
M403 436 75 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=46900 $D=1
M404 6 435 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=42270 $D=1
M405 7 436 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=46900 $D=1
M406 437 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=42270 $D=1
M407 438 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=46900 $D=1
M408 435 431 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=42270 $D=1
M409 436 432 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=46900 $D=1
M410 437 76 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=42270 $D=1
M411 438 76 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=46900 $D=1
M412 249 77 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=42270 $D=1
M413 250 77 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=46900 $D=1
M414 439 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=42270 $D=1
M415 440 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=46900 $D=1
M416 6 78 441 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=42270 $D=1
M417 7 78 442 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=46900 $D=1
M418 443 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=42270 $D=1
M419 444 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=46900 $D=1
M420 445 78 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=42270 $D=1
M421 446 78 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=46900 $D=1
M422 6 445 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=42270 $D=1
M423 7 446 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=46900 $D=1
M424 447 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=42270 $D=1
M425 448 751 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=46900 $D=1
M426 445 441 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=42270 $D=1
M427 446 442 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=46900 $D=1
M428 447 79 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=42270 $D=1
M429 448 79 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=46900 $D=1
M430 249 80 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=42270 $D=1
M431 250 80 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=46900 $D=1
M432 449 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=42270 $D=1
M433 450 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=46900 $D=1
M434 6 81 451 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=42270 $D=1
M435 7 81 452 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=46900 $D=1
M436 453 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=42270 $D=1
M437 454 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=46900 $D=1
M438 455 81 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=42270 $D=1
M439 456 81 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=46900 $D=1
M440 6 455 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=42270 $D=1
M441 7 456 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=46900 $D=1
M442 457 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=42270 $D=1
M443 458 753 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=46900 $D=1
M444 455 451 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=42270 $D=1
M445 456 452 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=46900 $D=1
M446 457 82 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=42270 $D=1
M447 458 82 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=46900 $D=1
M448 249 83 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=42270 $D=1
M449 250 83 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=46900 $D=1
M450 459 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=42270 $D=1
M451 460 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=46900 $D=1
M452 6 84 461 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=42270 $D=1
M453 7 84 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=46900 $D=1
M454 463 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=42270 $D=1
M455 464 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=46900 $D=1
M456 465 84 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=42270 $D=1
M457 466 84 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=46900 $D=1
M458 6 465 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=42270 $D=1
M459 7 466 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=46900 $D=1
M460 467 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=42270 $D=1
M461 468 755 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=46900 $D=1
M462 465 461 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=42270 $D=1
M463 466 462 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=46900 $D=1
M464 467 85 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=42270 $D=1
M465 468 85 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=46900 $D=1
M466 249 86 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=42270 $D=1
M467 250 86 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=46900 $D=1
M468 469 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=42270 $D=1
M469 470 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=46900 $D=1
M470 6 87 471 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=42270 $D=1
M471 7 87 472 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=46900 $D=1
M472 473 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=42270 $D=1
M473 474 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=46900 $D=1
M474 475 87 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=42270 $D=1
M475 476 87 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=46900 $D=1
M476 6 475 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=42270 $D=1
M477 7 476 757 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=46900 $D=1
M478 477 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=42270 $D=1
M479 478 757 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=46900 $D=1
M480 475 471 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=42270 $D=1
M481 476 472 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=46900 $D=1
M482 477 88 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=42270 $D=1
M483 478 88 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=46900 $D=1
M484 249 89 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=42270 $D=1
M485 250 89 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=46900 $D=1
M486 479 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=42270 $D=1
M487 480 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=46900 $D=1
M488 6 90 481 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=42270 $D=1
M489 7 90 482 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=46900 $D=1
M490 483 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=42270 $D=1
M491 484 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=46900 $D=1
M492 485 90 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=42270 $D=1
M493 486 90 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=46900 $D=1
M494 6 485 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=42270 $D=1
M495 7 486 759 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=46900 $D=1
M496 487 758 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=42270 $D=1
M497 488 759 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=46900 $D=1
M498 485 481 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=42270 $D=1
M499 486 482 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=46900 $D=1
M500 487 91 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=42270 $D=1
M501 488 91 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=46900 $D=1
M502 249 92 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=42270 $D=1
M503 250 92 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=46900 $D=1
M504 489 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=42270 $D=1
M505 490 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=46900 $D=1
M506 6 93 491 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=42270 $D=1
M507 7 93 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=46900 $D=1
M508 493 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=42270 $D=1
M509 494 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=46900 $D=1
M510 495 93 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=42270 $D=1
M511 496 93 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=46900 $D=1
M512 6 495 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=42270 $D=1
M513 7 496 761 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=46900 $D=1
M514 497 760 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=42270 $D=1
M515 498 761 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=46900 $D=1
M516 495 491 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=42270 $D=1
M517 496 492 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=46900 $D=1
M518 497 94 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=42270 $D=1
M519 498 94 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=46900 $D=1
M520 249 95 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=42270 $D=1
M521 250 95 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=46900 $D=1
M522 499 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=42270 $D=1
M523 500 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=46900 $D=1
M524 6 96 501 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=42270 $D=1
M525 7 96 502 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=46900 $D=1
M526 503 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=42270 $D=1
M527 504 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=46900 $D=1
M528 505 96 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=42270 $D=1
M529 506 96 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=46900 $D=1
M530 6 505 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=42270 $D=1
M531 7 506 763 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=46900 $D=1
M532 507 762 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=42270 $D=1
M533 508 763 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=46900 $D=1
M534 505 501 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=42270 $D=1
M535 506 502 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=46900 $D=1
M536 507 97 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=42270 $D=1
M537 508 97 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=46900 $D=1
M538 249 98 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=42270 $D=1
M539 250 98 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=46900 $D=1
M540 509 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=42270 $D=1
M541 510 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=46900 $D=1
M542 6 99 511 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=42270 $D=1
M543 7 99 512 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=46900 $D=1
M544 513 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=42270 $D=1
M545 514 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=46900 $D=1
M546 515 99 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=42270 $D=1
M547 516 99 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=46900 $D=1
M548 6 515 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=42270 $D=1
M549 7 516 765 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=46900 $D=1
M550 517 764 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=42270 $D=1
M551 518 765 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=46900 $D=1
M552 515 511 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=42270 $D=1
M553 516 512 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=46900 $D=1
M554 517 100 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=42270 $D=1
M555 518 100 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=46900 $D=1
M556 249 101 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=42270 $D=1
M557 250 101 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=46900 $D=1
M558 519 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=42270 $D=1
M559 520 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=46900 $D=1
M560 6 102 521 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=42270 $D=1
M561 7 102 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=46900 $D=1
M562 523 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=42270 $D=1
M563 524 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=46900 $D=1
M564 525 102 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=42270 $D=1
M565 526 102 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=46900 $D=1
M566 6 525 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=42270 $D=1
M567 7 526 767 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=46900 $D=1
M568 527 766 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=42270 $D=1
M569 528 767 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=46900 $D=1
M570 525 521 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=42270 $D=1
M571 526 522 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=46900 $D=1
M572 527 103 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=42270 $D=1
M573 528 103 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=46900 $D=1
M574 249 104 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=42270 $D=1
M575 250 104 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=46900 $D=1
M576 529 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=42270 $D=1
M577 530 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=46900 $D=1
M578 6 105 531 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=42270 $D=1
M579 7 105 532 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=46900 $D=1
M580 533 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=42270 $D=1
M581 534 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=46900 $D=1
M582 535 105 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=42270 $D=1
M583 536 105 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=46900 $D=1
M584 6 535 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=42270 $D=1
M585 7 536 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=46900 $D=1
M586 537 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=42270 $D=1
M587 538 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=46900 $D=1
M588 535 531 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=42270 $D=1
M589 536 532 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=46900 $D=1
M590 537 106 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=42270 $D=1
M591 538 106 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=46900 $D=1
M592 249 110 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=42270 $D=1
M593 250 110 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=46900 $D=1
M594 539 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=42270 $D=1
M595 540 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=46900 $D=1
M596 6 111 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=42270 $D=1
M597 7 111 542 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=46900 $D=1
M598 543 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=42270 $D=1
M599 544 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=46900 $D=1
M600 545 111 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=42270 $D=1
M601 546 111 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=46900 $D=1
M602 6 545 770 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=42270 $D=1
M603 7 546 771 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=46900 $D=1
M604 547 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=42270 $D=1
M605 548 771 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=46900 $D=1
M606 545 541 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=42270 $D=1
M607 546 542 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=46900 $D=1
M608 547 112 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=42270 $D=1
M609 548 112 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=46900 $D=1
M610 249 114 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=42270 $D=1
M611 250 114 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=46900 $D=1
M612 549 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=42270 $D=1
M613 550 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=46900 $D=1
M614 6 115 551 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=42270 $D=1
M615 7 115 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=46900 $D=1
M616 553 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=42270 $D=1
M617 554 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=46900 $D=1
M618 6 116 245 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=42270 $D=1
M619 7 116 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=46900 $D=1
M620 249 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=42270 $D=1
M621 250 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=46900 $D=1
M622 6 557 555 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=42270 $D=1
M623 7 558 556 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=46900 $D=1
M624 557 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=42270 $D=1
M625 558 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=46900 $D=1
M626 772 245 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=42270 $D=1
M627 773 246 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=46900 $D=1
M628 559 555 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=42270 $D=1
M629 560 556 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=46900 $D=1
M630 6 559 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=42270 $D=1
M631 7 560 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=46900 $D=1
M632 774 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=42270 $D=1
M633 775 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=46900 $D=1
M634 559 557 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=42270 $D=1
M635 560 558 775 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=46900 $D=1
M636 6 565 563 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=42270 $D=1
M637 7 566 564 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=46900 $D=1
M638 565 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=42270 $D=1
M639 566 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=46900 $D=1
M640 776 249 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=42270 $D=1
M641 777 250 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=46900 $D=1
M642 567 563 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=42270 $D=1
M643 568 564 777 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=46900 $D=1
M644 6 567 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=42270 $D=1
M645 7 568 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=46900 $D=1
M646 778 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=42270 $D=1
M647 779 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=46900 $D=1
M648 567 565 778 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=42270 $D=1
M649 568 566 779 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=46900 $D=1
M650 569 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=42270 $D=1
M651 570 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=46900 $D=1
M652 571 569 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=42270 $D=1
M653 572 570 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=46900 $D=1
M654 121 120 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=42270 $D=1
M655 122 120 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=46900 $D=1
M656 573 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=42270 $D=1
M657 574 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=46900 $D=1
M658 575 573 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=42270 $D=1
M659 576 574 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=46900 $D=1
M660 780 123 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=42270 $D=1
M661 781 123 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=46900 $D=1
M662 6 118 780 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=42270 $D=1
M663 7 119 781 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=46900 $D=1
M664 577 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=42270 $D=1
M665 578 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=46900 $D=1
M666 579 577 575 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=42270 $D=1
M667 580 578 576 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=46900 $D=1
M668 12 124 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=42270 $D=1
M669 13 124 580 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=46900 $D=1
M670 583 581 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=42270 $D=1
M671 584 582 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=46900 $D=1
M672 6 587 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=42270 $D=1
M673 7 588 586 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=46900 $D=1
M674 589 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=42270 $D=1
M675 590 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=46900 $D=1
M676 587 589 581 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=42270 $D=1
M677 588 590 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=46900 $D=1
M678 583 571 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=42270 $D=1
M679 584 572 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=46900 $D=1
M680 591 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=42270 $D=1
M681 592 586 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=46900 $D=1
M682 125 591 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=42270 $D=1
M683 581 592 580 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=46900 $D=1
M684 571 585 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=42270 $D=1
M685 572 586 581 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=46900 $D=1
M686 593 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=42270 $D=1
M687 594 581 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=46900 $D=1
M688 595 585 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=42270 $D=1
M689 596 586 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=46900 $D=1
M690 597 595 593 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=42270 $D=1
M691 598 596 594 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=46900 $D=1
M692 579 585 597 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=42270 $D=1
M693 580 586 598 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=46900 $D=1
M694 599 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=42270 $D=1
M695 600 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=46900 $D=1
M696 6 579 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=42270 $D=1
M697 7 580 600 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=46900 $D=1
M698 601 597 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=42270 $D=1
M699 602 598 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=46900 $D=1
M700 800 571 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=42270 $D=1
M701 801 572 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=46900 $D=1
M702 603 579 800 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=42270 $D=1
M703 604 580 801 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=46900 $D=1
M704 802 571 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=42270 $D=1
M705 803 572 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=46900 $D=1
M706 605 579 802 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=42270 $D=1
M707 606 580 803 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=46900 $D=1
M708 609 571 607 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=42270 $D=1
M709 610 572 608 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=46900 $D=1
M710 607 579 609 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=42270 $D=1
M711 608 580 610 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=46900 $D=1
M712 6 605 607 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=42270 $D=1
M713 7 606 608 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=46900 $D=1
M714 611 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=42270 $D=1
M715 612 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=46900 $D=1
M716 613 611 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=42270 $D=1
M717 614 612 600 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=46900 $D=1
M718 603 128 613 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=42270 $D=1
M719 604 128 614 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=46900 $D=1
M720 615 611 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=42270 $D=1
M721 616 612 602 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=46900 $D=1
M722 609 128 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=42270 $D=1
M723 610 128 616 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=46900 $D=1
M724 617 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=42270 $D=1
M725 618 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=46900 $D=1
M726 619 617 615 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=42270 $D=1
M727 620 618 616 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=46900 $D=1
M728 613 129 619 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=42270 $D=1
M729 614 129 620 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=46900 $D=1
M730 14 619 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=42270 $D=1
M731 15 620 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=46900 $D=1
M732 621 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=42270 $D=1
M733 622 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=46900 $D=1
M734 623 621 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=42270 $D=1
M735 624 622 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=46900 $D=1
M736 133 130 623 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=42270 $D=1
M737 134 130 624 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=46900 $D=1
M738 625 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=42270 $D=1
M739 626 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=46900 $D=1
M740 627 625 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=42270 $D=1
M741 628 626 136 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=46900 $D=1
M742 137 130 627 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=42270 $D=1
M743 138 130 628 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=46900 $D=1
M744 629 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=42270 $D=1
M745 630 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=46900 $D=1
M746 631 629 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=42270 $D=1
M747 632 630 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=46900 $D=1
M748 139 130 631 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=42270 $D=1
M749 109 130 632 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=46900 $D=1
M750 633 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=42270 $D=1
M751 634 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=46900 $D=1
M752 635 633 140 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=42270 $D=1
M753 636 634 141 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=46900 $D=1
M754 142 130 635 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=42270 $D=1
M755 143 130 636 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=46900 $D=1
M756 637 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=42270 $D=1
M757 638 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=46900 $D=1
M758 639 637 122 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=42270 $D=1
M759 640 638 144 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=46900 $D=1
M760 145 130 639 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=42270 $D=1
M761 145 130 640 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=46900 $D=1
M762 6 571 782 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=42270 $D=1
M763 7 572 783 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=46900 $D=1
M764 134 782 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=42270 $D=1
M765 131 783 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=46900 $D=1
M766 641 146 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=42270 $D=1
M767 642 146 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=46900 $D=1
M768 147 641 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=42270 $D=1
M769 148 642 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=46900 $D=1
M770 623 146 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=42270 $D=1
M771 624 146 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=46900 $D=1
M772 643 149 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=42270 $D=1
M773 644 149 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=46900 $D=1
M774 150 643 147 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=42270 $D=1
M775 107 644 148 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=46900 $D=1
M776 627 149 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=42270 $D=1
M777 628 149 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=46900 $D=1
M778 645 151 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=42270 $D=1
M779 646 151 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=46900 $D=1
M780 150 645 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=42270 $D=1
M781 107 646 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=46900 $D=1
M782 631 151 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=42270 $D=1
M783 632 151 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=46900 $D=1
M784 647 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=42270 $D=1
M785 648 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=46900 $D=1
M786 153 647 150 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=42270 $D=1
M787 154 648 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=46900 $D=1
M788 635 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=42270 $D=1
M789 636 152 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=46900 $D=1
M790 649 155 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=42270 $D=1
M791 650 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=46900 $D=1
M792 221 649 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=42270 $D=1
M793 222 650 154 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=46900 $D=1
M794 639 155 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=42270 $D=1
M795 640 155 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=46900 $D=1
M796 651 156 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=42270 $D=1
M797 652 156 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=46900 $D=1
M798 653 651 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=42270 $D=1
M799 654 652 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=46900 $D=1
M800 12 156 653 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=42270 $D=1
M801 13 156 654 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=46900 $D=1
M802 804 561 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=42270 $D=1
M803 805 562 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=46900 $D=1
M804 655 653 804 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=42270 $D=1
M805 656 654 805 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=46900 $D=1
M806 659 561 657 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=42270 $D=1
M807 660 562 658 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=46900 $D=1
M808 657 653 659 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=42270 $D=1
M809 658 654 660 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=46900 $D=1
M810 6 655 657 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=42270 $D=1
M811 7 656 658 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=46900 $D=1
M812 806 157 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=42270 $D=1
M813 807 661 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=46900 $D=1
M814 784 659 806 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=42270 $D=1
M815 785 660 807 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=46900 $D=1
M816 661 784 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=42270 $D=1
M817 158 785 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=46900 $D=1
M818 662 561 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=42270 $D=1
M819 663 562 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=46900 $D=1
M820 6 664 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=42270 $D=1
M821 7 665 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=46900 $D=1
M822 664 653 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=42270 $D=1
M823 665 654 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=46900 $D=1
M824 808 662 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=42270 $D=1
M825 809 663 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=46900 $D=1
M826 666 157 808 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=42270 $D=1
M827 667 661 809 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=46900 $D=1
M828 669 159 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=42270 $D=1
M829 670 668 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=46900 $D=1
M830 810 666 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=42270 $D=1
M831 811 667 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=46900 $D=1
M832 668 669 810 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=42270 $D=1
M833 160 670 811 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=46900 $D=1
M834 672 671 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=42270 $D=1
M835 673 161 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=46900 $D=1
M836 6 676 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=42270 $D=1
M837 7 677 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=46900 $D=1
M838 678 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=42270 $D=1
M839 679 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=46900 $D=1
M840 676 678 671 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=42270 $D=1
M841 677 679 161 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=46900 $D=1
M842 672 121 676 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=42270 $D=1
M843 673 122 677 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=46900 $D=1
M844 680 674 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=42270 $D=1
M845 681 675 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=46900 $D=1
M846 162 680 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=42270 $D=1
M847 671 681 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=46900 $D=1
M848 121 674 162 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=42270 $D=1
M849 122 675 671 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=46900 $D=1
M850 682 162 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=42270 $D=1
M851 683 671 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=46900 $D=1
M852 684 674 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=42270 $D=1
M853 685 675 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=46900 $D=1
M854 223 684 682 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=42270 $D=1
M855 224 685 683 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=46900 $D=1
M856 6 674 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=42270 $D=1
M857 7 675 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=46900 $D=1
M858 686 163 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=42270 $D=1
M859 687 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=46900 $D=1
M860 688 686 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=42270 $D=1
M861 689 687 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=46900 $D=1
M862 14 163 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=42270 $D=1
M863 15 163 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=46900 $D=1
M864 690 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=42270 $D=1
M865 691 164 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=46900 $D=1
M866 164 690 688 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=42270 $D=1
M867 164 691 689 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=46900 $D=1
M868 6 164 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=42270 $D=1
M869 7 164 164 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=46900 $D=1
M870 692 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=42270 $D=1
M871 693 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=46900 $D=1
M872 6 692 694 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=42270 $D=1
M873 7 693 695 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=46900 $D=1
M874 696 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=42270 $D=1
M875 697 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=46900 $D=1
M876 698 692 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=42270 $D=1
M877 699 693 164 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=46900 $D=1
M878 6 698 786 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=42270 $D=1
M879 7 699 787 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=46900 $D=1
M880 700 786 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=42270 $D=1
M881 701 787 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=46900 $D=1
M882 698 694 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=42270 $D=1
M883 699 695 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=46900 $D=1
M884 702 117 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=42270 $D=1
M885 703 117 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=46900 $D=1
M886 6 706 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=42270 $D=1
M887 7 707 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=46900 $D=1
M888 706 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=42270 $D=1
M889 707 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=46900 $D=1
M890 788 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=42270 $D=1
M891 789 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=46900 $D=1
M892 708 704 788 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=42270 $D=1
M893 709 705 789 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=46900 $D=1
M894 6 708 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=42270 $D=1
M895 7 709 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=46900 $D=1
M896 790 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=42270 $D=1
M897 791 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=46900 $D=1
M898 708 706 790 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=42270 $D=1
M899 709 707 791 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=46900 $D=1
M900 197 1 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=43520 $D=0
M901 198 1 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=48150 $D=0
M902 199 1 2 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=43520 $D=0
M903 200 1 3 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=48150 $D=0
M904 6 197 199 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=43520 $D=0
M905 7 198 200 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=48150 $D=0
M906 201 1 4 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=43520 $D=0
M907 202 1 4 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=48150 $D=0
M908 5 197 201 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=43520 $D=0
M909 5 198 202 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=48150 $D=0
M910 203 1 6 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=43520 $D=0
M911 204 1 7 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=48150 $D=0
M912 6 197 203 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=43520 $D=0
M913 7 198 204 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=48150 $D=0
M914 207 9 203 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=43520 $D=0
M915 208 9 204 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=48150 $D=0
M916 205 9 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=43520 $D=0
M917 206 9 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=48150 $D=0
M918 209 9 201 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=43520 $D=0
M919 210 9 202 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=48150 $D=0
M920 199 205 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=43520 $D=0
M921 200 206 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=48150 $D=0
M922 211 10 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=43520 $D=0
M923 212 10 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=48150 $D=0
M924 213 10 209 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=43520 $D=0
M925 214 10 210 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=48150 $D=0
M926 207 211 213 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=43520 $D=0
M927 208 212 214 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=48150 $D=0
M928 215 11 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=43520 $D=0
M929 216 11 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=48150 $D=0
M930 217 11 6 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=43520 $D=0
M931 218 11 7 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=48150 $D=0
M932 12 215 217 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=43520 $D=0
M933 13 216 218 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=48150 $D=0
M934 219 11 14 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=43520 $D=0
M935 220 11 15 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=48150 $D=0
M936 221 215 219 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=43520 $D=0
M937 222 216 220 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=48150 $D=0
M938 225 11 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=43520 $D=0
M939 226 11 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=48150 $D=0
M940 213 215 225 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=43520 $D=0
M941 214 216 226 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=48150 $D=0
M942 229 16 225 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=43520 $D=0
M943 230 16 226 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=48150 $D=0
M944 227 16 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=43520 $D=0
M945 228 16 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=48150 $D=0
M946 231 16 219 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=43520 $D=0
M947 232 16 220 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=48150 $D=0
M948 217 227 231 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=43520 $D=0
M949 218 228 232 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=48150 $D=0
M950 233 17 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=43520 $D=0
M951 234 17 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=48150 $D=0
M952 235 17 231 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=43520 $D=0
M953 236 17 232 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=48150 $D=0
M954 229 233 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=43520 $D=0
M955 230 234 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=48150 $D=0
M956 165 18 237 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=43520 $D=0
M957 166 18 238 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=48150 $D=0
M958 239 19 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=43520 $D=0
M959 240 19 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=48150 $D=0
M960 241 237 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=43520 $D=0
M961 242 238 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=48150 $D=0
M962 165 241 710 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=43520 $D=0
M963 166 242 711 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=48150 $D=0
M964 243 710 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=43520 $D=0
M965 244 711 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=48150 $D=0
M966 241 18 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=43520 $D=0
M967 242 18 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=48150 $D=0
M968 243 239 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=43520 $D=0
M969 244 240 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=48150 $D=0
M970 249 247 243 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=43520 $D=0
M971 250 248 244 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=48150 $D=0
M972 247 20 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=43520 $D=0
M973 248 20 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=48150 $D=0
M974 165 21 251 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=43520 $D=0
M975 166 21 252 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=48150 $D=0
M976 253 22 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=43520 $D=0
M977 254 22 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=48150 $D=0
M978 255 251 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=43520 $D=0
M979 256 252 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=48150 $D=0
M980 165 255 712 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=43520 $D=0
M981 166 256 713 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=48150 $D=0
M982 257 712 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=43520 $D=0
M983 258 713 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=48150 $D=0
M984 255 21 257 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=43520 $D=0
M985 256 21 258 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=48150 $D=0
M986 257 253 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=43520 $D=0
M987 258 254 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=48150 $D=0
M988 249 259 257 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=43520 $D=0
M989 250 260 258 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=48150 $D=0
M990 259 23 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=43520 $D=0
M991 260 23 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=48150 $D=0
M992 165 24 261 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=43520 $D=0
M993 166 24 262 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=48150 $D=0
M994 263 25 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=43520 $D=0
M995 264 25 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=48150 $D=0
M996 265 261 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=43520 $D=0
M997 266 262 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=48150 $D=0
M998 165 265 714 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=43520 $D=0
M999 166 266 715 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=48150 $D=0
M1000 267 714 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=43520 $D=0
M1001 268 715 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=48150 $D=0
M1002 265 24 267 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=43520 $D=0
M1003 266 24 268 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=48150 $D=0
M1004 267 263 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=43520 $D=0
M1005 268 264 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=48150 $D=0
M1006 249 269 267 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=43520 $D=0
M1007 250 270 268 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=48150 $D=0
M1008 269 26 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=43520 $D=0
M1009 270 26 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=48150 $D=0
M1010 165 27 271 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=43520 $D=0
M1011 166 27 272 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=48150 $D=0
M1012 273 28 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=43520 $D=0
M1013 274 28 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=48150 $D=0
M1014 275 271 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=43520 $D=0
M1015 276 272 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=48150 $D=0
M1016 165 275 716 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=43520 $D=0
M1017 166 276 717 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=48150 $D=0
M1018 277 716 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=43520 $D=0
M1019 278 717 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=48150 $D=0
M1020 275 27 277 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=43520 $D=0
M1021 276 27 278 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=48150 $D=0
M1022 277 273 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=43520 $D=0
M1023 278 274 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=48150 $D=0
M1024 249 279 277 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=43520 $D=0
M1025 250 280 278 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=48150 $D=0
M1026 279 29 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=43520 $D=0
M1027 280 29 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=48150 $D=0
M1028 165 30 281 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=43520 $D=0
M1029 166 30 282 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=48150 $D=0
M1030 283 31 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=43520 $D=0
M1031 284 31 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=48150 $D=0
M1032 285 281 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=43520 $D=0
M1033 286 282 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=48150 $D=0
M1034 165 285 718 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=43520 $D=0
M1035 166 286 719 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=48150 $D=0
M1036 287 718 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=43520 $D=0
M1037 288 719 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=48150 $D=0
M1038 285 30 287 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=43520 $D=0
M1039 286 30 288 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=48150 $D=0
M1040 287 283 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=43520 $D=0
M1041 288 284 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=48150 $D=0
M1042 249 289 287 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=43520 $D=0
M1043 250 290 288 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=48150 $D=0
M1044 289 32 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=43520 $D=0
M1045 290 32 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=48150 $D=0
M1046 165 33 291 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=43520 $D=0
M1047 166 33 292 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=48150 $D=0
M1048 293 34 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=43520 $D=0
M1049 294 34 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=48150 $D=0
M1050 295 291 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=43520 $D=0
M1051 296 292 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=48150 $D=0
M1052 165 295 720 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=43520 $D=0
M1053 166 296 721 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=48150 $D=0
M1054 297 720 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=43520 $D=0
M1055 298 721 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=48150 $D=0
M1056 295 33 297 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=43520 $D=0
M1057 296 33 298 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=48150 $D=0
M1058 297 293 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=43520 $D=0
M1059 298 294 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=48150 $D=0
M1060 249 299 297 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=43520 $D=0
M1061 250 300 298 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=48150 $D=0
M1062 299 35 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=43520 $D=0
M1063 300 35 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=48150 $D=0
M1064 165 36 301 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=43520 $D=0
M1065 166 36 302 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=48150 $D=0
M1066 303 37 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=43520 $D=0
M1067 304 37 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=48150 $D=0
M1068 305 301 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=43520 $D=0
M1069 306 302 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=48150 $D=0
M1070 165 305 722 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=43520 $D=0
M1071 166 306 723 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=48150 $D=0
M1072 307 722 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=43520 $D=0
M1073 308 723 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=48150 $D=0
M1074 305 36 307 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=43520 $D=0
M1075 306 36 308 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=48150 $D=0
M1076 307 303 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=43520 $D=0
M1077 308 304 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=48150 $D=0
M1078 249 309 307 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=43520 $D=0
M1079 250 310 308 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=48150 $D=0
M1080 309 38 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=43520 $D=0
M1081 310 38 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=48150 $D=0
M1082 165 39 311 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=43520 $D=0
M1083 166 39 312 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=48150 $D=0
M1084 313 40 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=43520 $D=0
M1085 314 40 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=48150 $D=0
M1086 315 311 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=43520 $D=0
M1087 316 312 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=48150 $D=0
M1088 165 315 724 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=43520 $D=0
M1089 166 316 725 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=48150 $D=0
M1090 317 724 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=43520 $D=0
M1091 318 725 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=48150 $D=0
M1092 315 39 317 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=43520 $D=0
M1093 316 39 318 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=48150 $D=0
M1094 317 313 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=43520 $D=0
M1095 318 314 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=48150 $D=0
M1096 249 319 317 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=43520 $D=0
M1097 250 320 318 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=48150 $D=0
M1098 319 41 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=43520 $D=0
M1099 320 41 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=48150 $D=0
M1100 165 42 321 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=43520 $D=0
M1101 166 42 322 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=48150 $D=0
M1102 323 43 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=43520 $D=0
M1103 324 43 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=48150 $D=0
M1104 325 321 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=43520 $D=0
M1105 326 322 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=48150 $D=0
M1106 165 325 726 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=43520 $D=0
M1107 166 326 727 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=48150 $D=0
M1108 327 726 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=43520 $D=0
M1109 328 727 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=48150 $D=0
M1110 325 42 327 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=43520 $D=0
M1111 326 42 328 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=48150 $D=0
M1112 327 323 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=43520 $D=0
M1113 328 324 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=48150 $D=0
M1114 249 329 327 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=43520 $D=0
M1115 250 330 328 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=48150 $D=0
M1116 329 44 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=43520 $D=0
M1117 330 44 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=48150 $D=0
M1118 165 45 331 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=43520 $D=0
M1119 166 45 332 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=48150 $D=0
M1120 333 46 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=43520 $D=0
M1121 334 46 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=48150 $D=0
M1122 335 331 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=43520 $D=0
M1123 336 332 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=48150 $D=0
M1124 165 335 728 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=43520 $D=0
M1125 166 336 729 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=48150 $D=0
M1126 337 728 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=43520 $D=0
M1127 338 729 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=48150 $D=0
M1128 335 45 337 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=43520 $D=0
M1129 336 45 338 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=48150 $D=0
M1130 337 333 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=43520 $D=0
M1131 338 334 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=48150 $D=0
M1132 249 339 337 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=43520 $D=0
M1133 250 340 338 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=48150 $D=0
M1134 339 47 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=43520 $D=0
M1135 340 47 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=48150 $D=0
M1136 165 48 341 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=43520 $D=0
M1137 166 48 342 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=48150 $D=0
M1138 343 49 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=43520 $D=0
M1139 344 49 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=48150 $D=0
M1140 345 341 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=43520 $D=0
M1141 346 342 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=48150 $D=0
M1142 165 345 730 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=43520 $D=0
M1143 166 346 731 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=48150 $D=0
M1144 347 730 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=43520 $D=0
M1145 348 731 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=48150 $D=0
M1146 345 48 347 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=43520 $D=0
M1147 346 48 348 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=48150 $D=0
M1148 347 343 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=43520 $D=0
M1149 348 344 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=48150 $D=0
M1150 249 349 347 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=43520 $D=0
M1151 250 350 348 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=48150 $D=0
M1152 349 50 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=43520 $D=0
M1153 350 50 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=48150 $D=0
M1154 165 51 351 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=43520 $D=0
M1155 166 51 352 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=48150 $D=0
M1156 353 52 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=43520 $D=0
M1157 354 52 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=48150 $D=0
M1158 355 351 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=43520 $D=0
M1159 356 352 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=48150 $D=0
M1160 165 355 732 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=43520 $D=0
M1161 166 356 733 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=48150 $D=0
M1162 357 732 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=43520 $D=0
M1163 358 733 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=48150 $D=0
M1164 355 51 357 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=43520 $D=0
M1165 356 51 358 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=48150 $D=0
M1166 357 353 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=43520 $D=0
M1167 358 354 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=48150 $D=0
M1168 249 359 357 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=43520 $D=0
M1169 250 360 358 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=48150 $D=0
M1170 359 53 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=43520 $D=0
M1171 360 53 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=48150 $D=0
M1172 165 54 361 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=43520 $D=0
M1173 166 54 362 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=48150 $D=0
M1174 363 55 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=43520 $D=0
M1175 364 55 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=48150 $D=0
M1176 365 361 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=43520 $D=0
M1177 366 362 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=48150 $D=0
M1178 165 365 734 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=43520 $D=0
M1179 166 366 735 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=48150 $D=0
M1180 367 734 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=43520 $D=0
M1181 368 735 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=48150 $D=0
M1182 365 54 367 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=43520 $D=0
M1183 366 54 368 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=48150 $D=0
M1184 367 363 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=43520 $D=0
M1185 368 364 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=48150 $D=0
M1186 249 369 367 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=43520 $D=0
M1187 250 370 368 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=48150 $D=0
M1188 369 56 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=43520 $D=0
M1189 370 56 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=48150 $D=0
M1190 165 57 371 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=43520 $D=0
M1191 166 57 372 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=48150 $D=0
M1192 373 58 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=43520 $D=0
M1193 374 58 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=48150 $D=0
M1194 375 371 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=43520 $D=0
M1195 376 372 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=48150 $D=0
M1196 165 375 736 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=43520 $D=0
M1197 166 376 737 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=48150 $D=0
M1198 377 736 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=43520 $D=0
M1199 378 737 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=48150 $D=0
M1200 375 57 377 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=43520 $D=0
M1201 376 57 378 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=48150 $D=0
M1202 377 373 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=43520 $D=0
M1203 378 374 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=48150 $D=0
M1204 249 379 377 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=43520 $D=0
M1205 250 380 378 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=48150 $D=0
M1206 379 59 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=43520 $D=0
M1207 380 59 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=48150 $D=0
M1208 165 60 381 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=43520 $D=0
M1209 166 60 382 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=48150 $D=0
M1210 383 61 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=43520 $D=0
M1211 384 61 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=48150 $D=0
M1212 385 381 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=43520 $D=0
M1213 386 382 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=48150 $D=0
M1214 165 385 738 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=43520 $D=0
M1215 166 386 739 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=48150 $D=0
M1216 387 738 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=43520 $D=0
M1217 388 739 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=48150 $D=0
M1218 385 60 387 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=43520 $D=0
M1219 386 60 388 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=48150 $D=0
M1220 387 383 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=43520 $D=0
M1221 388 384 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=48150 $D=0
M1222 249 389 387 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=43520 $D=0
M1223 250 390 388 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=48150 $D=0
M1224 389 62 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=43520 $D=0
M1225 390 62 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=48150 $D=0
M1226 165 63 391 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=43520 $D=0
M1227 166 63 392 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=48150 $D=0
M1228 393 64 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=43520 $D=0
M1229 394 64 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=48150 $D=0
M1230 395 391 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=43520 $D=0
M1231 396 392 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=48150 $D=0
M1232 165 395 740 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=43520 $D=0
M1233 166 396 741 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=48150 $D=0
M1234 397 740 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=43520 $D=0
M1235 398 741 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=48150 $D=0
M1236 395 63 397 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=43520 $D=0
M1237 396 63 398 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=48150 $D=0
M1238 397 393 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=43520 $D=0
M1239 398 394 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=48150 $D=0
M1240 249 399 397 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=43520 $D=0
M1241 250 400 398 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=48150 $D=0
M1242 399 65 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=43520 $D=0
M1243 400 65 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=48150 $D=0
M1244 165 66 401 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=43520 $D=0
M1245 166 66 402 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=48150 $D=0
M1246 403 67 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=43520 $D=0
M1247 404 67 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=48150 $D=0
M1248 405 401 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=43520 $D=0
M1249 406 402 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=48150 $D=0
M1250 165 405 742 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=43520 $D=0
M1251 166 406 743 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=48150 $D=0
M1252 407 742 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=43520 $D=0
M1253 408 743 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=48150 $D=0
M1254 405 66 407 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=43520 $D=0
M1255 406 66 408 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=48150 $D=0
M1256 407 403 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=43520 $D=0
M1257 408 404 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=48150 $D=0
M1258 249 409 407 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=43520 $D=0
M1259 250 410 408 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=48150 $D=0
M1260 409 68 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=43520 $D=0
M1261 410 68 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=48150 $D=0
M1262 165 69 411 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=43520 $D=0
M1263 166 69 412 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=48150 $D=0
M1264 413 70 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=43520 $D=0
M1265 414 70 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=48150 $D=0
M1266 415 411 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=43520 $D=0
M1267 416 412 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=48150 $D=0
M1268 165 415 744 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=43520 $D=0
M1269 166 416 745 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=48150 $D=0
M1270 417 744 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=43520 $D=0
M1271 418 745 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=48150 $D=0
M1272 415 69 417 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=43520 $D=0
M1273 416 69 418 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=48150 $D=0
M1274 417 413 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=43520 $D=0
M1275 418 414 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=48150 $D=0
M1276 249 419 417 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=43520 $D=0
M1277 250 420 418 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=48150 $D=0
M1278 419 71 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=43520 $D=0
M1279 420 71 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=48150 $D=0
M1280 165 72 421 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=43520 $D=0
M1281 166 72 422 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=48150 $D=0
M1282 423 73 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=43520 $D=0
M1283 424 73 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=48150 $D=0
M1284 425 421 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=43520 $D=0
M1285 426 422 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=48150 $D=0
M1286 165 425 746 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=43520 $D=0
M1287 166 426 747 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=48150 $D=0
M1288 427 746 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=43520 $D=0
M1289 428 747 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=48150 $D=0
M1290 425 72 427 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=43520 $D=0
M1291 426 72 428 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=48150 $D=0
M1292 427 423 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=43520 $D=0
M1293 428 424 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=48150 $D=0
M1294 249 429 427 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=43520 $D=0
M1295 250 430 428 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=48150 $D=0
M1296 429 74 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=43520 $D=0
M1297 430 74 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=48150 $D=0
M1298 165 75 431 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=43520 $D=0
M1299 166 75 432 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=48150 $D=0
M1300 433 76 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=43520 $D=0
M1301 434 76 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=48150 $D=0
M1302 435 431 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=43520 $D=0
M1303 436 432 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=48150 $D=0
M1304 165 435 748 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=43520 $D=0
M1305 166 436 749 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=48150 $D=0
M1306 437 748 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=43520 $D=0
M1307 438 749 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=48150 $D=0
M1308 435 75 437 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=43520 $D=0
M1309 436 75 438 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=48150 $D=0
M1310 437 433 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=43520 $D=0
M1311 438 434 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=48150 $D=0
M1312 249 439 437 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=43520 $D=0
M1313 250 440 438 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=48150 $D=0
M1314 439 77 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=43520 $D=0
M1315 440 77 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=48150 $D=0
M1316 165 78 441 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=43520 $D=0
M1317 166 78 442 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=48150 $D=0
M1318 443 79 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=43520 $D=0
M1319 444 79 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=48150 $D=0
M1320 445 441 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=43520 $D=0
M1321 446 442 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=48150 $D=0
M1322 165 445 750 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=43520 $D=0
M1323 166 446 751 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=48150 $D=0
M1324 447 750 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=43520 $D=0
M1325 448 751 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=48150 $D=0
M1326 445 78 447 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=43520 $D=0
M1327 446 78 448 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=48150 $D=0
M1328 447 443 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=43520 $D=0
M1329 448 444 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=48150 $D=0
M1330 249 449 447 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=43520 $D=0
M1331 250 450 448 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=48150 $D=0
M1332 449 80 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=43520 $D=0
M1333 450 80 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=48150 $D=0
M1334 165 81 451 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=43520 $D=0
M1335 166 81 452 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=48150 $D=0
M1336 453 82 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=43520 $D=0
M1337 454 82 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=48150 $D=0
M1338 455 451 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=43520 $D=0
M1339 456 452 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=48150 $D=0
M1340 165 455 752 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=43520 $D=0
M1341 166 456 753 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=48150 $D=0
M1342 457 752 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=43520 $D=0
M1343 458 753 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=48150 $D=0
M1344 455 81 457 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=43520 $D=0
M1345 456 81 458 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=48150 $D=0
M1346 457 453 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=43520 $D=0
M1347 458 454 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=48150 $D=0
M1348 249 459 457 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=43520 $D=0
M1349 250 460 458 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=48150 $D=0
M1350 459 83 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=43520 $D=0
M1351 460 83 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=48150 $D=0
M1352 165 84 461 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=43520 $D=0
M1353 166 84 462 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=48150 $D=0
M1354 463 85 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=43520 $D=0
M1355 464 85 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=48150 $D=0
M1356 465 461 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=43520 $D=0
M1357 466 462 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=48150 $D=0
M1358 165 465 754 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=43520 $D=0
M1359 166 466 755 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=48150 $D=0
M1360 467 754 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=43520 $D=0
M1361 468 755 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=48150 $D=0
M1362 465 84 467 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=43520 $D=0
M1363 466 84 468 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=48150 $D=0
M1364 467 463 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=43520 $D=0
M1365 468 464 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=48150 $D=0
M1366 249 469 467 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=43520 $D=0
M1367 250 470 468 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=48150 $D=0
M1368 469 86 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=43520 $D=0
M1369 470 86 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=48150 $D=0
M1370 165 87 471 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=43520 $D=0
M1371 166 87 472 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=48150 $D=0
M1372 473 88 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=43520 $D=0
M1373 474 88 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=48150 $D=0
M1374 475 471 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=43520 $D=0
M1375 476 472 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=48150 $D=0
M1376 165 475 756 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=43520 $D=0
M1377 166 476 757 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=48150 $D=0
M1378 477 756 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=43520 $D=0
M1379 478 757 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=48150 $D=0
M1380 475 87 477 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=43520 $D=0
M1381 476 87 478 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=48150 $D=0
M1382 477 473 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=43520 $D=0
M1383 478 474 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=48150 $D=0
M1384 249 479 477 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=43520 $D=0
M1385 250 480 478 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=48150 $D=0
M1386 479 89 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=43520 $D=0
M1387 480 89 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=48150 $D=0
M1388 165 90 481 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=43520 $D=0
M1389 166 90 482 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=48150 $D=0
M1390 483 91 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=43520 $D=0
M1391 484 91 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=48150 $D=0
M1392 485 481 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=43520 $D=0
M1393 486 482 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=48150 $D=0
M1394 165 485 758 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=43520 $D=0
M1395 166 486 759 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=48150 $D=0
M1396 487 758 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=43520 $D=0
M1397 488 759 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=48150 $D=0
M1398 485 90 487 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=43520 $D=0
M1399 486 90 488 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=48150 $D=0
M1400 487 483 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=43520 $D=0
M1401 488 484 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=48150 $D=0
M1402 249 489 487 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=43520 $D=0
M1403 250 490 488 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=48150 $D=0
M1404 489 92 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=43520 $D=0
M1405 490 92 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=48150 $D=0
M1406 165 93 491 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=43520 $D=0
M1407 166 93 492 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=48150 $D=0
M1408 493 94 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=43520 $D=0
M1409 494 94 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=48150 $D=0
M1410 495 491 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=43520 $D=0
M1411 496 492 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=48150 $D=0
M1412 165 495 760 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=43520 $D=0
M1413 166 496 761 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=48150 $D=0
M1414 497 760 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=43520 $D=0
M1415 498 761 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=48150 $D=0
M1416 495 93 497 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=43520 $D=0
M1417 496 93 498 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=48150 $D=0
M1418 497 493 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=43520 $D=0
M1419 498 494 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=48150 $D=0
M1420 249 499 497 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=43520 $D=0
M1421 250 500 498 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=48150 $D=0
M1422 499 95 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=43520 $D=0
M1423 500 95 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=48150 $D=0
M1424 165 96 501 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=43520 $D=0
M1425 166 96 502 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=48150 $D=0
M1426 503 97 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=43520 $D=0
M1427 504 97 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=48150 $D=0
M1428 505 501 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=43520 $D=0
M1429 506 502 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=48150 $D=0
M1430 165 505 762 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=43520 $D=0
M1431 166 506 763 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=48150 $D=0
M1432 507 762 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=43520 $D=0
M1433 508 763 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=48150 $D=0
M1434 505 96 507 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=43520 $D=0
M1435 506 96 508 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=48150 $D=0
M1436 507 503 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=43520 $D=0
M1437 508 504 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=48150 $D=0
M1438 249 509 507 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=43520 $D=0
M1439 250 510 508 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=48150 $D=0
M1440 509 98 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=43520 $D=0
M1441 510 98 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=48150 $D=0
M1442 165 99 511 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=43520 $D=0
M1443 166 99 512 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=48150 $D=0
M1444 513 100 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=43520 $D=0
M1445 514 100 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=48150 $D=0
M1446 515 511 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=43520 $D=0
M1447 516 512 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=48150 $D=0
M1448 165 515 764 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=43520 $D=0
M1449 166 516 765 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=48150 $D=0
M1450 517 764 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=43520 $D=0
M1451 518 765 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=48150 $D=0
M1452 515 99 517 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=43520 $D=0
M1453 516 99 518 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=48150 $D=0
M1454 517 513 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=43520 $D=0
M1455 518 514 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=48150 $D=0
M1456 249 519 517 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=43520 $D=0
M1457 250 520 518 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=48150 $D=0
M1458 519 101 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=43520 $D=0
M1459 520 101 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=48150 $D=0
M1460 165 102 521 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=43520 $D=0
M1461 166 102 522 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=48150 $D=0
M1462 523 103 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=43520 $D=0
M1463 524 103 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=48150 $D=0
M1464 525 521 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=43520 $D=0
M1465 526 522 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=48150 $D=0
M1466 165 525 766 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=43520 $D=0
M1467 166 526 767 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=48150 $D=0
M1468 527 766 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=43520 $D=0
M1469 528 767 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=48150 $D=0
M1470 525 102 527 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=43520 $D=0
M1471 526 102 528 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=48150 $D=0
M1472 527 523 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=43520 $D=0
M1473 528 524 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=48150 $D=0
M1474 249 529 527 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=43520 $D=0
M1475 250 530 528 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=48150 $D=0
M1476 529 104 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=43520 $D=0
M1477 530 104 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=48150 $D=0
M1478 165 105 531 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=43520 $D=0
M1479 166 105 532 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=48150 $D=0
M1480 533 106 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=43520 $D=0
M1481 534 106 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=48150 $D=0
M1482 535 531 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=43520 $D=0
M1483 536 532 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=48150 $D=0
M1484 165 535 768 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=43520 $D=0
M1485 166 536 769 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=48150 $D=0
M1486 537 768 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=43520 $D=0
M1487 538 769 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=48150 $D=0
M1488 535 105 537 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=43520 $D=0
M1489 536 105 538 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=48150 $D=0
M1490 537 533 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=43520 $D=0
M1491 538 534 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=48150 $D=0
M1492 249 539 537 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=43520 $D=0
M1493 250 540 538 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=48150 $D=0
M1494 539 110 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=43520 $D=0
M1495 540 110 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=48150 $D=0
M1496 165 111 541 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=43520 $D=0
M1497 166 111 542 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=48150 $D=0
M1498 543 112 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=43520 $D=0
M1499 544 112 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=48150 $D=0
M1500 545 541 235 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=43520 $D=0
M1501 546 542 236 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=48150 $D=0
M1502 165 545 770 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=43520 $D=0
M1503 166 546 771 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=48150 $D=0
M1504 547 770 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=43520 $D=0
M1505 548 771 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=48150 $D=0
M1506 545 111 547 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=43520 $D=0
M1507 546 111 548 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=48150 $D=0
M1508 547 543 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=43520 $D=0
M1509 548 544 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=48150 $D=0
M1510 249 549 547 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=43520 $D=0
M1511 250 550 548 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=48150 $D=0
M1512 549 114 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=43520 $D=0
M1513 550 114 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=48150 $D=0
M1514 165 115 551 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=43520 $D=0
M1515 166 115 552 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=48150 $D=0
M1516 553 116 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=43520 $D=0
M1517 554 116 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=48150 $D=0
M1518 6 553 245 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=43520 $D=0
M1519 7 554 246 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=48150 $D=0
M1520 249 551 6 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=43520 $D=0
M1521 250 552 7 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=48150 $D=0
M1522 165 557 555 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=43520 $D=0
M1523 166 558 556 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=48150 $D=0
M1524 557 117 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=43520 $D=0
M1525 558 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=48150 $D=0
M1526 772 245 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=43520 $D=0
M1527 773 246 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=48150 $D=0
M1528 559 557 772 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=43520 $D=0
M1529 560 558 773 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=48150 $D=0
M1530 165 559 561 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=43520 $D=0
M1531 166 560 562 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=48150 $D=0
M1532 774 561 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=43520 $D=0
M1533 775 562 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=48150 $D=0
M1534 559 555 774 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=43520 $D=0
M1535 560 556 775 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=48150 $D=0
M1536 165 565 563 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=43520 $D=0
M1537 166 566 564 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=48150 $D=0
M1538 565 117 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=43520 $D=0
M1539 566 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=48150 $D=0
M1540 776 249 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=43520 $D=0
M1541 777 250 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=48150 $D=0
M1542 567 565 776 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=43520 $D=0
M1543 568 566 777 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=48150 $D=0
M1544 165 567 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=43520 $D=0
M1545 166 568 119 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=48150 $D=0
M1546 778 118 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=43520 $D=0
M1547 779 119 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=48150 $D=0
M1548 567 563 778 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=43520 $D=0
M1549 568 564 779 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=48150 $D=0
M1550 569 120 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=43520 $D=0
M1551 570 120 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=48150 $D=0
M1552 571 120 561 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=43520 $D=0
M1553 572 120 562 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=48150 $D=0
M1554 121 569 571 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=43520 $D=0
M1555 122 570 572 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=48150 $D=0
M1556 573 123 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=43520 $D=0
M1557 574 123 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=48150 $D=0
M1558 575 123 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=43520 $D=0
M1559 576 123 119 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=48150 $D=0
M1560 780 573 575 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=43520 $D=0
M1561 781 574 576 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=48150 $D=0
M1562 165 118 780 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=43520 $D=0
M1563 166 119 781 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=48150 $D=0
M1564 577 124 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=43520 $D=0
M1565 578 124 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=48150 $D=0
M1566 579 124 575 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=43520 $D=0
M1567 580 124 576 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=48150 $D=0
M1568 12 577 579 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=43520 $D=0
M1569 13 578 580 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=48150 $D=0
M1570 583 581 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=43520 $D=0
M1571 584 582 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=48150 $D=0
M1572 165 587 585 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=43520 $D=0
M1573 166 588 586 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=48150 $D=0
M1574 589 571 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=43520 $D=0
M1575 590 572 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=48150 $D=0
M1576 587 571 581 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=43520 $D=0
M1577 588 572 582 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=48150 $D=0
M1578 583 589 587 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=43520 $D=0
M1579 584 590 588 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=48150 $D=0
M1580 591 585 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=43520 $D=0
M1581 592 586 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=48150 $D=0
M1582 125 585 579 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=43520 $D=0
M1583 581 586 580 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=48150 $D=0
M1584 571 591 125 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=43520 $D=0
M1585 572 592 581 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=48150 $D=0
M1586 593 125 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=43520 $D=0
M1587 594 581 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=48150 $D=0
M1588 595 585 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=43520 $D=0
M1589 596 586 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=48150 $D=0
M1590 597 585 593 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=43520 $D=0
M1591 598 586 594 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=48150 $D=0
M1592 579 595 597 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=43520 $D=0
M1593 580 596 598 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=48150 $D=0
M1594 792 571 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=43160 $D=0
M1595 793 572 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=47790 $D=0
M1596 599 579 792 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=43160 $D=0
M1597 600 580 793 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=47790 $D=0
M1598 601 597 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=43520 $D=0
M1599 602 598 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=48150 $D=0
M1600 603 571 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=43520 $D=0
M1601 604 572 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=48150 $D=0
M1602 165 579 603 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=43520 $D=0
M1603 166 580 604 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=48150 $D=0
M1604 605 571 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=43520 $D=0
M1605 606 572 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=48150 $D=0
M1606 165 579 605 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=43520 $D=0
M1607 166 580 606 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=48150 $D=0
M1608 794 571 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=43340 $D=0
M1609 795 572 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=47970 $D=0
M1610 609 579 794 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=43340 $D=0
M1611 610 580 795 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=47970 $D=0
M1612 165 605 609 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=43520 $D=0
M1613 166 606 610 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=48150 $D=0
M1614 611 128 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=43520 $D=0
M1615 612 128 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=48150 $D=0
M1616 613 128 599 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=43520 $D=0
M1617 614 128 600 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=48150 $D=0
M1618 603 611 613 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=43520 $D=0
M1619 604 612 614 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=48150 $D=0
M1620 615 128 601 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=43520 $D=0
M1621 616 128 602 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=48150 $D=0
M1622 609 611 615 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=43520 $D=0
M1623 610 612 616 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=48150 $D=0
M1624 617 129 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=43520 $D=0
M1625 618 129 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=48150 $D=0
M1626 619 129 615 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=43520 $D=0
M1627 620 129 616 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=48150 $D=0
M1628 613 617 619 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=43520 $D=0
M1629 614 618 620 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=48150 $D=0
M1630 14 619 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=43520 $D=0
M1631 15 620 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=48150 $D=0
M1632 621 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=43520 $D=0
M1633 622 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=48150 $D=0
M1634 623 130 131 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=43520 $D=0
M1635 624 130 132 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=48150 $D=0
M1636 133 621 623 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=43520 $D=0
M1637 134 622 624 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=48150 $D=0
M1638 625 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=43520 $D=0
M1639 626 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=48150 $D=0
M1640 627 130 135 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=43520 $D=0
M1641 628 130 136 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=48150 $D=0
M1642 137 625 627 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=43520 $D=0
M1643 138 626 628 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=48150 $D=0
M1644 629 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=43520 $D=0
M1645 630 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=48150 $D=0
M1646 631 130 127 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=43520 $D=0
M1647 632 130 126 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=48150 $D=0
M1648 139 629 631 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=43520 $D=0
M1649 109 630 632 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=48150 $D=0
M1650 633 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=43520 $D=0
M1651 634 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=48150 $D=0
M1652 635 130 140 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=43520 $D=0
M1653 636 130 141 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=48150 $D=0
M1654 142 633 635 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=43520 $D=0
M1655 143 634 636 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=48150 $D=0
M1656 637 130 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=43520 $D=0
M1657 638 130 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=48150 $D=0
M1658 639 130 122 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=43520 $D=0
M1659 640 130 144 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=48150 $D=0
M1660 145 637 639 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=43520 $D=0
M1661 145 638 640 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=48150 $D=0
M1662 165 571 782 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=43520 $D=0
M1663 166 572 783 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=48150 $D=0
M1664 134 782 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=43520 $D=0
M1665 131 783 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=48150 $D=0
M1666 641 146 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=43520 $D=0
M1667 642 146 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=48150 $D=0
M1668 147 146 134 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=43520 $D=0
M1669 148 146 131 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=48150 $D=0
M1670 623 641 147 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=43520 $D=0
M1671 624 642 148 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=48150 $D=0
M1672 643 149 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=43520 $D=0
M1673 644 149 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=48150 $D=0
M1674 150 149 147 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=43520 $D=0
M1675 107 149 148 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=48150 $D=0
M1676 627 643 150 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=43520 $D=0
M1677 628 644 107 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=48150 $D=0
M1678 645 151 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=43520 $D=0
M1679 646 151 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=48150 $D=0
M1680 150 151 150 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=43520 $D=0
M1681 107 151 107 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=48150 $D=0
M1682 631 645 150 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=43520 $D=0
M1683 632 646 107 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=48150 $D=0
M1684 647 152 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=43520 $D=0
M1685 648 152 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=48150 $D=0
M1686 153 152 150 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=43520 $D=0
M1687 154 152 107 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=48150 $D=0
M1688 635 647 153 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=43520 $D=0
M1689 636 648 154 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=48150 $D=0
M1690 649 155 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=43520 $D=0
M1691 650 155 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=48150 $D=0
M1692 221 155 153 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=43520 $D=0
M1693 222 155 154 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=48150 $D=0
M1694 639 649 221 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=43520 $D=0
M1695 640 650 222 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=48150 $D=0
M1696 651 156 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=43520 $D=0
M1697 652 156 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=48150 $D=0
M1698 653 156 118 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=43520 $D=0
M1699 654 156 119 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=48150 $D=0
M1700 12 651 653 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=43520 $D=0
M1701 13 652 654 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=48150 $D=0
M1702 655 561 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=43520 $D=0
M1703 656 562 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=48150 $D=0
M1704 165 653 655 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=43520 $D=0
M1705 166 654 656 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=48150 $D=0
M1706 796 561 165 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=43340 $D=0
M1707 797 562 166 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=47970 $D=0
M1708 659 653 796 165 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=43340 $D=0
M1709 660 654 797 166 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=47970 $D=0
M1710 165 655 659 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=43520 $D=0
M1711 166 656 660 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=48150 $D=0
M1712 784 157 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=43520 $D=0
M1713 785 661 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=48150 $D=0
M1714 165 659 784 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=43520 $D=0
M1715 166 660 785 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=48150 $D=0
M1716 661 784 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=43520 $D=0
M1717 158 785 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=48150 $D=0
M1718 798 561 165 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=43160 $D=0
M1719 799 562 166 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=47790 $D=0
M1720 662 664 798 165 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=43160 $D=0
M1721 663 665 799 166 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=47790 $D=0
M1722 664 653 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=43520 $D=0
M1723 665 654 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=48150 $D=0
M1724 666 662 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=43520 $D=0
M1725 667 663 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=48150 $D=0
M1726 165 157 666 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=43520 $D=0
M1727 166 661 667 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=48150 $D=0
M1728 669 159 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=43520 $D=0
M1729 670 668 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=48150 $D=0
M1730 668 666 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=43520 $D=0
M1731 160 667 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=48150 $D=0
M1732 165 669 668 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=43520 $D=0
M1733 166 670 160 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=48150 $D=0
M1734 672 671 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=43520 $D=0
M1735 673 161 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=48150 $D=0
M1736 165 676 674 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=43520 $D=0
M1737 166 677 675 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=48150 $D=0
M1738 678 121 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=43520 $D=0
M1739 679 122 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=48150 $D=0
M1740 676 121 671 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=43520 $D=0
M1741 677 122 161 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=48150 $D=0
M1742 672 678 676 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=43520 $D=0
M1743 673 679 677 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=48150 $D=0
M1744 680 674 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=43520 $D=0
M1745 681 675 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=48150 $D=0
M1746 162 674 6 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=43520 $D=0
M1747 671 675 7 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=48150 $D=0
M1748 121 680 162 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=43520 $D=0
M1749 122 681 671 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=48150 $D=0
M1750 682 162 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=43520 $D=0
M1751 683 671 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=48150 $D=0
M1752 684 674 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=43520 $D=0
M1753 685 675 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=48150 $D=0
M1754 223 674 682 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=43520 $D=0
M1755 224 675 683 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=48150 $D=0
M1756 6 684 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=43520 $D=0
M1757 7 685 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=48150 $D=0
M1758 686 163 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=43520 $D=0
M1759 687 163 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=48150 $D=0
M1760 688 163 223 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=43520 $D=0
M1761 689 163 224 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=48150 $D=0
M1762 14 686 688 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=43520 $D=0
M1763 15 687 689 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=48150 $D=0
M1764 690 164 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=43520 $D=0
M1765 691 164 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=48150 $D=0
M1766 164 164 688 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=43520 $D=0
M1767 164 164 689 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=48150 $D=0
M1768 6 690 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=43520 $D=0
M1769 7 691 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=48150 $D=0
M1770 692 117 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=43520 $D=0
M1771 693 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=48150 $D=0
M1772 165 692 694 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=43520 $D=0
M1773 166 693 695 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=48150 $D=0
M1774 696 117 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=43520 $D=0
M1775 697 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=48150 $D=0
M1776 698 694 164 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=43520 $D=0
M1777 699 695 164 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=48150 $D=0
M1778 165 698 786 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=43520 $D=0
M1779 166 699 787 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=48150 $D=0
M1780 700 786 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=43520 $D=0
M1781 701 787 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=48150 $D=0
M1782 698 692 700 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=43520 $D=0
M1783 699 693 701 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=48150 $D=0
M1784 702 696 700 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=43520 $D=0
M1785 703 697 701 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=48150 $D=0
M1786 165 706 704 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=43520 $D=0
M1787 166 707 705 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=48150 $D=0
M1788 706 117 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=43520 $D=0
M1789 707 117 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=48150 $D=0
M1790 788 702 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=43520 $D=0
M1791 789 703 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=48150 $D=0
M1792 708 706 788 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=43520 $D=0
M1793 709 707 789 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=48150 $D=0
M1794 165 708 121 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=43520 $D=0
M1795 166 709 122 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=48150 $D=0
M1796 790 121 165 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=43520 $D=0
M1797 791 122 166 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=48150 $D=0
M1798 708 704 790 165 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=43520 $D=0
M1799 709 705 791 166 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=48150 $D=0
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 109 110 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168
** N=808 EP=165 IP=1514 FDC=1800
M0 195 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=33010 $D=1
M1 196 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=37640 $D=1
M2 197 195 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=33010 $D=1
M3 198 196 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=37640 $D=1
M4 6 1 197 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=33010 $D=1
M5 7 1 198 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=37640 $D=1
M6 199 195 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=33010 $D=1
M7 200 196 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=37640 $D=1
M8 5 1 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=33010 $D=1
M9 5 1 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=37640 $D=1
M10 201 195 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=33010 $D=1
M11 202 196 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=37640 $D=1
M12 6 1 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=33010 $D=1
M13 7 1 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=37640 $D=1
M14 205 203 201 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=33010 $D=1
M15 206 204 202 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=37640 $D=1
M16 203 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=33010 $D=1
M17 204 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=37640 $D=1
M18 207 203 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=33010 $D=1
M19 208 204 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=37640 $D=1
M20 197 9 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=33010 $D=1
M21 198 9 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=37640 $D=1
M22 209 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=33010 $D=1
M23 210 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=37640 $D=1
M24 211 209 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=33010 $D=1
M25 212 210 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=37640 $D=1
M26 205 10 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=33010 $D=1
M27 206 10 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=37640 $D=1
M28 213 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=33010 $D=1
M29 214 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=37640 $D=1
M30 215 213 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=33010 $D=1
M31 216 214 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=37640 $D=1
M32 12 11 215 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=33010 $D=1
M33 13 11 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=37640 $D=1
M34 217 213 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=33010 $D=1
M35 218 214 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=37640 $D=1
M36 219 11 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=33010 $D=1
M37 220 11 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=37640 $D=1
M38 223 213 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=33010 $D=1
M39 224 214 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=37640 $D=1
M40 211 11 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=33010 $D=1
M41 212 11 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=37640 $D=1
M42 227 225 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=33010 $D=1
M43 228 226 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=37640 $D=1
M44 225 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=33010 $D=1
M45 226 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=37640 $D=1
M46 229 225 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=33010 $D=1
M47 230 226 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=37640 $D=1
M48 215 16 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=33010 $D=1
M49 216 16 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=37640 $D=1
M50 231 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=33010 $D=1
M51 232 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=37640 $D=1
M52 233 231 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=33010 $D=1
M53 234 232 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=37640 $D=1
M54 227 17 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=33010 $D=1
M55 228 17 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=37640 $D=1
M56 6 18 235 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=33010 $D=1
M57 7 18 236 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=37640 $D=1
M58 237 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=33010 $D=1
M59 238 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=37640 $D=1
M60 239 18 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=33010 $D=1
M61 240 18 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=37640 $D=1
M62 6 239 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=33010 $D=1
M63 7 240 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=37640 $D=1
M64 241 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=33010 $D=1
M65 242 708 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=37640 $D=1
M66 239 235 241 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=33010 $D=1
M67 240 236 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=37640 $D=1
M68 241 19 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=33010 $D=1
M69 242 19 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=37640 $D=1
M70 247 20 241 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=33010 $D=1
M71 248 20 242 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=37640 $D=1
M72 245 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=33010 $D=1
M73 246 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=37640 $D=1
M74 6 21 249 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=33010 $D=1
M75 7 21 250 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=37640 $D=1
M76 251 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=33010 $D=1
M77 252 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=37640 $D=1
M78 253 21 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=33010 $D=1
M79 254 21 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=37640 $D=1
M80 6 253 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=33010 $D=1
M81 7 254 710 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=37640 $D=1
M82 255 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=33010 $D=1
M83 256 710 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=37640 $D=1
M84 253 249 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=33010 $D=1
M85 254 250 256 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=37640 $D=1
M86 255 22 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=33010 $D=1
M87 256 22 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=37640 $D=1
M88 247 23 255 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=33010 $D=1
M89 248 23 256 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=37640 $D=1
M90 257 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=33010 $D=1
M91 258 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=37640 $D=1
M92 6 24 259 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=33010 $D=1
M93 7 24 260 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=37640 $D=1
M94 261 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=33010 $D=1
M95 262 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=37640 $D=1
M96 263 24 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=33010 $D=1
M97 264 24 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=37640 $D=1
M98 6 263 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=33010 $D=1
M99 7 264 712 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=37640 $D=1
M100 265 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=33010 $D=1
M101 266 712 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=37640 $D=1
M102 263 259 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=33010 $D=1
M103 264 260 266 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=37640 $D=1
M104 265 25 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=33010 $D=1
M105 266 25 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=37640 $D=1
M106 247 26 265 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=33010 $D=1
M107 248 26 266 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=37640 $D=1
M108 267 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=33010 $D=1
M109 268 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=37640 $D=1
M110 6 27 269 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=33010 $D=1
M111 7 27 270 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=37640 $D=1
M112 271 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=33010 $D=1
M113 272 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=37640 $D=1
M114 273 27 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=33010 $D=1
M115 274 27 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=37640 $D=1
M116 6 273 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=33010 $D=1
M117 7 274 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=37640 $D=1
M118 275 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=33010 $D=1
M119 276 714 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=37640 $D=1
M120 273 269 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=33010 $D=1
M121 274 270 276 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=37640 $D=1
M122 275 28 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=33010 $D=1
M123 276 28 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=37640 $D=1
M124 247 29 275 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=33010 $D=1
M125 248 29 276 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=37640 $D=1
M126 277 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=33010 $D=1
M127 278 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=37640 $D=1
M128 6 30 279 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=33010 $D=1
M129 7 30 280 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=37640 $D=1
M130 281 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=33010 $D=1
M131 282 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=37640 $D=1
M132 283 30 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=33010 $D=1
M133 284 30 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=37640 $D=1
M134 6 283 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=33010 $D=1
M135 7 284 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=37640 $D=1
M136 285 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=33010 $D=1
M137 286 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=37640 $D=1
M138 283 279 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=33010 $D=1
M139 284 280 286 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=37640 $D=1
M140 285 31 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=33010 $D=1
M141 286 31 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=37640 $D=1
M142 247 32 285 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=33010 $D=1
M143 248 32 286 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=37640 $D=1
M144 287 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=33010 $D=1
M145 288 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=37640 $D=1
M146 6 33 289 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=33010 $D=1
M147 7 33 290 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=37640 $D=1
M148 291 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=33010 $D=1
M149 292 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=37640 $D=1
M150 293 33 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=33010 $D=1
M151 294 33 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=37640 $D=1
M152 6 293 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=33010 $D=1
M153 7 294 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=37640 $D=1
M154 295 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=33010 $D=1
M155 296 718 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=37640 $D=1
M156 293 289 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=33010 $D=1
M157 294 290 296 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=37640 $D=1
M158 295 34 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=33010 $D=1
M159 296 34 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=37640 $D=1
M160 247 35 295 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=33010 $D=1
M161 248 35 296 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=37640 $D=1
M162 297 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=33010 $D=1
M163 298 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=37640 $D=1
M164 6 36 299 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=33010 $D=1
M165 7 36 300 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=37640 $D=1
M166 301 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=33010 $D=1
M167 302 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=37640 $D=1
M168 303 36 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=33010 $D=1
M169 304 36 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=37640 $D=1
M170 6 303 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=33010 $D=1
M171 7 304 720 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=37640 $D=1
M172 305 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=33010 $D=1
M173 306 720 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=37640 $D=1
M174 303 299 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=33010 $D=1
M175 304 300 306 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=37640 $D=1
M176 305 37 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=33010 $D=1
M177 306 37 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=37640 $D=1
M178 247 38 305 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=33010 $D=1
M179 248 38 306 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=37640 $D=1
M180 307 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=33010 $D=1
M181 308 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=37640 $D=1
M182 6 39 309 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=33010 $D=1
M183 7 39 310 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=37640 $D=1
M184 311 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=33010 $D=1
M185 312 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=37640 $D=1
M186 313 39 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=33010 $D=1
M187 314 39 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=37640 $D=1
M188 6 313 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=33010 $D=1
M189 7 314 722 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=37640 $D=1
M190 315 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=33010 $D=1
M191 316 722 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=37640 $D=1
M192 313 309 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=33010 $D=1
M193 314 310 316 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=37640 $D=1
M194 315 40 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=33010 $D=1
M195 316 40 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=37640 $D=1
M196 247 41 315 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=33010 $D=1
M197 248 41 316 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=37640 $D=1
M198 317 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=33010 $D=1
M199 318 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=37640 $D=1
M200 6 42 319 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=33010 $D=1
M201 7 42 320 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=37640 $D=1
M202 321 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=33010 $D=1
M203 322 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=37640 $D=1
M204 323 42 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=33010 $D=1
M205 324 42 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=37640 $D=1
M206 6 323 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=33010 $D=1
M207 7 324 724 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=37640 $D=1
M208 325 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=33010 $D=1
M209 326 724 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=37640 $D=1
M210 323 319 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=33010 $D=1
M211 324 320 326 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=37640 $D=1
M212 325 43 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=33010 $D=1
M213 326 43 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=37640 $D=1
M214 247 44 325 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=33010 $D=1
M215 248 44 326 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=37640 $D=1
M216 327 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=33010 $D=1
M217 328 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=37640 $D=1
M218 6 45 329 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=33010 $D=1
M219 7 45 330 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=37640 $D=1
M220 331 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=33010 $D=1
M221 332 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=37640 $D=1
M222 333 45 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=33010 $D=1
M223 334 45 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=37640 $D=1
M224 6 333 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=33010 $D=1
M225 7 334 726 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=37640 $D=1
M226 335 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=33010 $D=1
M227 336 726 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=37640 $D=1
M228 333 329 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=33010 $D=1
M229 334 330 336 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=37640 $D=1
M230 335 46 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=33010 $D=1
M231 336 46 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=37640 $D=1
M232 247 47 335 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=33010 $D=1
M233 248 47 336 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=37640 $D=1
M234 337 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=33010 $D=1
M235 338 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=37640 $D=1
M236 6 48 339 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=33010 $D=1
M237 7 48 340 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=37640 $D=1
M238 341 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=33010 $D=1
M239 342 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=37640 $D=1
M240 343 48 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=33010 $D=1
M241 344 48 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=37640 $D=1
M242 6 343 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=33010 $D=1
M243 7 344 728 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=37640 $D=1
M244 345 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=33010 $D=1
M245 346 728 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=37640 $D=1
M246 343 339 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=33010 $D=1
M247 344 340 346 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=37640 $D=1
M248 345 49 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=33010 $D=1
M249 346 49 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=37640 $D=1
M250 247 50 345 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=33010 $D=1
M251 248 50 346 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=37640 $D=1
M252 347 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=33010 $D=1
M253 348 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=37640 $D=1
M254 6 51 349 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=33010 $D=1
M255 7 51 350 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=37640 $D=1
M256 351 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=33010 $D=1
M257 352 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=37640 $D=1
M258 353 51 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=33010 $D=1
M259 354 51 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=37640 $D=1
M260 6 353 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=33010 $D=1
M261 7 354 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=37640 $D=1
M262 355 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=33010 $D=1
M263 356 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=37640 $D=1
M264 353 349 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=33010 $D=1
M265 354 350 356 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=37640 $D=1
M266 355 52 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=33010 $D=1
M267 356 52 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=37640 $D=1
M268 247 53 355 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=33010 $D=1
M269 248 53 356 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=37640 $D=1
M270 357 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=33010 $D=1
M271 358 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=37640 $D=1
M272 6 54 359 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=33010 $D=1
M273 7 54 360 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=37640 $D=1
M274 361 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=33010 $D=1
M275 362 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=37640 $D=1
M276 363 54 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=33010 $D=1
M277 364 54 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=37640 $D=1
M278 6 363 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=33010 $D=1
M279 7 364 732 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=37640 $D=1
M280 365 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=33010 $D=1
M281 366 732 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=37640 $D=1
M282 363 359 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=33010 $D=1
M283 364 360 366 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=37640 $D=1
M284 365 55 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=33010 $D=1
M285 366 55 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=37640 $D=1
M286 247 56 365 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=33010 $D=1
M287 248 56 366 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=37640 $D=1
M288 367 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=33010 $D=1
M289 368 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=37640 $D=1
M290 6 57 369 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=33010 $D=1
M291 7 57 370 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=37640 $D=1
M292 371 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=33010 $D=1
M293 372 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=37640 $D=1
M294 373 57 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=33010 $D=1
M295 374 57 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=37640 $D=1
M296 6 373 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=33010 $D=1
M297 7 374 734 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=37640 $D=1
M298 375 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=33010 $D=1
M299 376 734 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=37640 $D=1
M300 373 369 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=33010 $D=1
M301 374 370 376 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=37640 $D=1
M302 375 58 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=33010 $D=1
M303 376 58 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=37640 $D=1
M304 247 59 375 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=33010 $D=1
M305 248 59 376 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=37640 $D=1
M306 377 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=33010 $D=1
M307 378 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=37640 $D=1
M308 6 60 379 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=33010 $D=1
M309 7 60 380 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=37640 $D=1
M310 381 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=33010 $D=1
M311 382 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=37640 $D=1
M312 383 60 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=33010 $D=1
M313 384 60 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=37640 $D=1
M314 6 383 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=33010 $D=1
M315 7 384 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=37640 $D=1
M316 385 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=33010 $D=1
M317 386 736 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=37640 $D=1
M318 383 379 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=33010 $D=1
M319 384 380 386 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=37640 $D=1
M320 385 61 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=33010 $D=1
M321 386 61 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=37640 $D=1
M322 247 62 385 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=33010 $D=1
M323 248 62 386 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=37640 $D=1
M324 387 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=33010 $D=1
M325 388 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=37640 $D=1
M326 6 63 389 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=33010 $D=1
M327 7 63 390 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=37640 $D=1
M328 391 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=33010 $D=1
M329 392 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=37640 $D=1
M330 393 63 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=33010 $D=1
M331 394 63 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=37640 $D=1
M332 6 393 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=33010 $D=1
M333 7 394 738 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=37640 $D=1
M334 395 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=33010 $D=1
M335 396 738 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=37640 $D=1
M336 393 389 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=33010 $D=1
M337 394 390 396 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=37640 $D=1
M338 395 64 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=33010 $D=1
M339 396 64 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=37640 $D=1
M340 247 65 395 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=33010 $D=1
M341 248 65 396 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=37640 $D=1
M342 397 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=33010 $D=1
M343 398 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=37640 $D=1
M344 6 66 399 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=33010 $D=1
M345 7 66 400 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=37640 $D=1
M346 401 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=33010 $D=1
M347 402 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=37640 $D=1
M348 403 66 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=33010 $D=1
M349 404 66 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=37640 $D=1
M350 6 403 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=33010 $D=1
M351 7 404 740 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=37640 $D=1
M352 405 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=33010 $D=1
M353 406 740 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=37640 $D=1
M354 403 399 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=33010 $D=1
M355 404 400 406 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=37640 $D=1
M356 405 67 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=33010 $D=1
M357 406 67 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=37640 $D=1
M358 247 68 405 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=33010 $D=1
M359 248 68 406 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=37640 $D=1
M360 407 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=33010 $D=1
M361 408 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=37640 $D=1
M362 6 69 409 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=33010 $D=1
M363 7 69 410 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=37640 $D=1
M364 411 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=33010 $D=1
M365 412 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=37640 $D=1
M366 413 69 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=33010 $D=1
M367 414 69 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=37640 $D=1
M368 6 413 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=33010 $D=1
M369 7 414 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=37640 $D=1
M370 415 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=33010 $D=1
M371 416 742 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=37640 $D=1
M372 413 409 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=33010 $D=1
M373 414 410 416 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=37640 $D=1
M374 415 70 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=33010 $D=1
M375 416 70 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=37640 $D=1
M376 247 71 415 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=33010 $D=1
M377 248 71 416 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=37640 $D=1
M378 417 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=33010 $D=1
M379 418 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=37640 $D=1
M380 6 72 419 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=33010 $D=1
M381 7 72 420 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=37640 $D=1
M382 421 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=33010 $D=1
M383 422 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=37640 $D=1
M384 423 72 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=33010 $D=1
M385 424 72 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=37640 $D=1
M386 6 423 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=33010 $D=1
M387 7 424 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=37640 $D=1
M388 425 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=33010 $D=1
M389 426 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=37640 $D=1
M390 423 419 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=33010 $D=1
M391 424 420 426 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=37640 $D=1
M392 425 73 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=33010 $D=1
M393 426 73 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=37640 $D=1
M394 247 74 425 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=33010 $D=1
M395 248 74 426 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=37640 $D=1
M396 427 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=33010 $D=1
M397 428 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=37640 $D=1
M398 6 75 429 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=33010 $D=1
M399 7 75 430 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=37640 $D=1
M400 431 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=33010 $D=1
M401 432 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=37640 $D=1
M402 433 75 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=33010 $D=1
M403 434 75 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=37640 $D=1
M404 6 433 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=33010 $D=1
M405 7 434 746 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=37640 $D=1
M406 435 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=33010 $D=1
M407 436 746 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=37640 $D=1
M408 433 429 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=33010 $D=1
M409 434 430 436 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=37640 $D=1
M410 435 76 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=33010 $D=1
M411 436 76 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=37640 $D=1
M412 247 77 435 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=33010 $D=1
M413 248 77 436 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=37640 $D=1
M414 437 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=33010 $D=1
M415 438 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=37640 $D=1
M416 6 78 439 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=33010 $D=1
M417 7 78 440 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=37640 $D=1
M418 441 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=33010 $D=1
M419 442 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=37640 $D=1
M420 443 78 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=33010 $D=1
M421 444 78 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=37640 $D=1
M422 6 443 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=33010 $D=1
M423 7 444 748 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=37640 $D=1
M424 445 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=33010 $D=1
M425 446 748 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=37640 $D=1
M426 443 439 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=33010 $D=1
M427 444 440 446 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=37640 $D=1
M428 445 79 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=33010 $D=1
M429 446 79 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=37640 $D=1
M430 247 80 445 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=33010 $D=1
M431 248 80 446 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=37640 $D=1
M432 447 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=33010 $D=1
M433 448 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=37640 $D=1
M434 6 81 449 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=33010 $D=1
M435 7 81 450 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=37640 $D=1
M436 451 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=33010 $D=1
M437 452 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=37640 $D=1
M438 453 81 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=33010 $D=1
M439 454 81 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=37640 $D=1
M440 6 453 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=33010 $D=1
M441 7 454 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=37640 $D=1
M442 455 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=33010 $D=1
M443 456 750 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=37640 $D=1
M444 453 449 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=33010 $D=1
M445 454 450 456 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=37640 $D=1
M446 455 82 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=33010 $D=1
M447 456 82 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=37640 $D=1
M448 247 83 455 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=33010 $D=1
M449 248 83 456 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=37640 $D=1
M450 457 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=33010 $D=1
M451 458 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=37640 $D=1
M452 6 84 459 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=33010 $D=1
M453 7 84 460 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=37640 $D=1
M454 461 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=33010 $D=1
M455 462 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=37640 $D=1
M456 463 84 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=33010 $D=1
M457 464 84 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=37640 $D=1
M458 6 463 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=33010 $D=1
M459 7 464 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=37640 $D=1
M460 465 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=33010 $D=1
M461 466 752 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=37640 $D=1
M462 463 459 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=33010 $D=1
M463 464 460 466 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=37640 $D=1
M464 465 85 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=33010 $D=1
M465 466 85 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=37640 $D=1
M466 247 86 465 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=33010 $D=1
M467 248 86 466 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=37640 $D=1
M468 467 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=33010 $D=1
M469 468 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=37640 $D=1
M470 6 87 469 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=33010 $D=1
M471 7 87 470 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=37640 $D=1
M472 471 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=33010 $D=1
M473 472 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=37640 $D=1
M474 473 87 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=33010 $D=1
M475 474 87 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=37640 $D=1
M476 6 473 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=33010 $D=1
M477 7 474 754 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=37640 $D=1
M478 475 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=33010 $D=1
M479 476 754 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=37640 $D=1
M480 473 469 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=33010 $D=1
M481 474 470 476 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=37640 $D=1
M482 475 88 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=33010 $D=1
M483 476 88 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=37640 $D=1
M484 247 89 475 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=33010 $D=1
M485 248 89 476 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=37640 $D=1
M486 477 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=33010 $D=1
M487 478 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=37640 $D=1
M488 6 90 479 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=33010 $D=1
M489 7 90 480 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=37640 $D=1
M490 481 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=33010 $D=1
M491 482 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=37640 $D=1
M492 483 90 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=33010 $D=1
M493 484 90 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=37640 $D=1
M494 6 483 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=33010 $D=1
M495 7 484 756 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=37640 $D=1
M496 485 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=33010 $D=1
M497 486 756 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=37640 $D=1
M498 483 479 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=33010 $D=1
M499 484 480 486 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=37640 $D=1
M500 485 91 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=33010 $D=1
M501 486 91 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=37640 $D=1
M502 247 92 485 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=33010 $D=1
M503 248 92 486 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=37640 $D=1
M504 487 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=33010 $D=1
M505 488 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=37640 $D=1
M506 6 93 489 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=33010 $D=1
M507 7 93 490 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=37640 $D=1
M508 491 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=33010 $D=1
M509 492 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=37640 $D=1
M510 493 93 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=33010 $D=1
M511 494 93 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=37640 $D=1
M512 6 493 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=33010 $D=1
M513 7 494 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=37640 $D=1
M514 495 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=33010 $D=1
M515 496 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=37640 $D=1
M516 493 489 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=33010 $D=1
M517 494 490 496 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=37640 $D=1
M518 495 94 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=33010 $D=1
M519 496 94 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=37640 $D=1
M520 247 95 495 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=33010 $D=1
M521 248 95 496 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=37640 $D=1
M522 497 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=33010 $D=1
M523 498 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=37640 $D=1
M524 6 96 499 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=33010 $D=1
M525 7 96 500 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=37640 $D=1
M526 501 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=33010 $D=1
M527 502 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=37640 $D=1
M528 503 96 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=33010 $D=1
M529 504 96 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=37640 $D=1
M530 6 503 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=33010 $D=1
M531 7 504 760 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=37640 $D=1
M532 505 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=33010 $D=1
M533 506 760 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=37640 $D=1
M534 503 499 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=33010 $D=1
M535 504 500 506 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=37640 $D=1
M536 505 97 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=33010 $D=1
M537 506 97 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=37640 $D=1
M538 247 98 505 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=33010 $D=1
M539 248 98 506 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=37640 $D=1
M540 507 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=33010 $D=1
M541 508 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=37640 $D=1
M542 6 99 509 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=33010 $D=1
M543 7 99 510 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=37640 $D=1
M544 511 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=33010 $D=1
M545 512 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=37640 $D=1
M546 513 99 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=33010 $D=1
M547 514 99 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=37640 $D=1
M548 6 513 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=33010 $D=1
M549 7 514 762 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=37640 $D=1
M550 515 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=33010 $D=1
M551 516 762 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=37640 $D=1
M552 513 509 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=33010 $D=1
M553 514 510 516 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=37640 $D=1
M554 515 100 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=33010 $D=1
M555 516 100 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=37640 $D=1
M556 247 101 515 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=33010 $D=1
M557 248 101 516 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=37640 $D=1
M558 517 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=33010 $D=1
M559 518 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=37640 $D=1
M560 6 102 519 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=33010 $D=1
M561 7 102 520 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=37640 $D=1
M562 521 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=33010 $D=1
M563 522 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=37640 $D=1
M564 523 102 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=33010 $D=1
M565 524 102 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=37640 $D=1
M566 6 523 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=33010 $D=1
M567 7 524 764 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=37640 $D=1
M568 525 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=33010 $D=1
M569 526 764 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=37640 $D=1
M570 523 519 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=33010 $D=1
M571 524 520 526 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=37640 $D=1
M572 525 103 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=33010 $D=1
M573 526 103 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=37640 $D=1
M574 247 104 525 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=33010 $D=1
M575 248 104 526 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=37640 $D=1
M576 527 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=33010 $D=1
M577 528 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=37640 $D=1
M578 6 105 529 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=33010 $D=1
M579 7 105 530 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=37640 $D=1
M580 531 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=33010 $D=1
M581 532 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=37640 $D=1
M582 533 105 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=33010 $D=1
M583 534 105 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=37640 $D=1
M584 6 533 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=33010 $D=1
M585 7 534 766 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=37640 $D=1
M586 535 765 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=33010 $D=1
M587 536 766 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=37640 $D=1
M588 533 529 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=33010 $D=1
M589 534 530 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=37640 $D=1
M590 535 106 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=33010 $D=1
M591 536 106 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=37640 $D=1
M592 247 110 535 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=33010 $D=1
M593 248 110 536 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=37640 $D=1
M594 537 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=33010 $D=1
M595 538 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=37640 $D=1
M596 6 112 539 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=33010 $D=1
M597 7 112 540 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=37640 $D=1
M598 541 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=33010 $D=1
M599 542 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=37640 $D=1
M600 543 112 233 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=33010 $D=1
M601 544 112 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=37640 $D=1
M602 6 543 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=33010 $D=1
M603 7 544 768 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=37640 $D=1
M604 545 767 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=33010 $D=1
M605 546 768 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=37640 $D=1
M606 543 539 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=33010 $D=1
M607 544 540 546 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=37640 $D=1
M608 545 113 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=33010 $D=1
M609 546 113 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=37640 $D=1
M610 247 114 545 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=33010 $D=1
M611 248 114 546 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=37640 $D=1
M612 547 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=33010 $D=1
M613 548 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=37640 $D=1
M614 6 115 549 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=33010 $D=1
M615 7 115 550 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=37640 $D=1
M616 551 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=33010 $D=1
M617 552 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=37640 $D=1
M618 6 116 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=33010 $D=1
M619 7 116 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=37640 $D=1
M620 247 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=33010 $D=1
M621 248 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=37640 $D=1
M622 6 555 553 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=33010 $D=1
M623 7 556 554 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=37640 $D=1
M624 555 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=33010 $D=1
M625 556 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=37640 $D=1
M626 769 243 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=33010 $D=1
M627 770 244 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=37640 $D=1
M628 557 553 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=33010 $D=1
M629 558 554 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=37640 $D=1
M630 6 557 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=33010 $D=1
M631 7 558 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=37640 $D=1
M632 771 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=33010 $D=1
M633 772 560 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=37640 $D=1
M634 557 555 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=33010 $D=1
M635 558 556 772 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=37640 $D=1
M636 6 563 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=33010 $D=1
M637 7 564 562 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=37640 $D=1
M638 563 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=33010 $D=1
M639 564 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=37640 $D=1
M640 773 247 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=33010 $D=1
M641 774 248 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=37640 $D=1
M642 565 561 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=33010 $D=1
M643 566 562 774 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=37640 $D=1
M644 6 565 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=33010 $D=1
M645 7 566 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=37640 $D=1
M646 775 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=33010 $D=1
M647 776 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=37640 $D=1
M648 565 563 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=33010 $D=1
M649 566 564 776 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=37640 $D=1
M650 567 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=33010 $D=1
M651 568 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=37640 $D=1
M652 569 567 559 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=33010 $D=1
M653 570 568 560 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=37640 $D=1
M654 121 120 569 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=33010 $D=1
M655 122 120 570 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=37640 $D=1
M656 571 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=33010 $D=1
M657 572 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=37640 $D=1
M658 573 571 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=33010 $D=1
M659 574 572 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=37640 $D=1
M660 777 123 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=33010 $D=1
M661 778 123 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=37640 $D=1
M662 6 118 777 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=33010 $D=1
M663 7 119 778 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=37640 $D=1
M664 575 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=33010 $D=1
M665 576 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=37640 $D=1
M666 577 575 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=33010 $D=1
M667 578 576 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=37640 $D=1
M668 12 124 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=33010 $D=1
M669 13 124 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=37640 $D=1
M670 580 579 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=33010 $D=1
M671 581 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=37640 $D=1
M672 6 584 582 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=33010 $D=1
M673 7 585 583 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=37640 $D=1
M674 586 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=33010 $D=1
M675 587 570 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=37640 $D=1
M676 584 586 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=33010 $D=1
M677 585 587 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=37640 $D=1
M678 580 569 584 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=33010 $D=1
M679 581 570 585 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=37640 $D=1
M680 588 582 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=33010 $D=1
M681 589 583 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=37640 $D=1
M682 126 588 577 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=33010 $D=1
M683 579 589 578 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=37640 $D=1
M684 569 582 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=33010 $D=1
M685 570 583 579 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=37640 $D=1
M686 590 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=33010 $D=1
M687 591 579 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=37640 $D=1
M688 592 582 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=33010 $D=1
M689 593 583 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=37640 $D=1
M690 594 592 590 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=33010 $D=1
M691 595 593 591 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=37640 $D=1
M692 577 582 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=33010 $D=1
M693 578 583 595 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=37640 $D=1
M694 596 569 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=33010 $D=1
M695 597 570 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=37640 $D=1
M696 6 577 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=33010 $D=1
M697 7 578 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=37640 $D=1
M698 598 594 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=33010 $D=1
M699 599 595 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=37640 $D=1
M700 797 569 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=33010 $D=1
M701 798 570 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=37640 $D=1
M702 600 577 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=33010 $D=1
M703 601 578 798 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=37640 $D=1
M704 799 569 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=33010 $D=1
M705 800 570 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=37640 $D=1
M706 602 577 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=33010 $D=1
M707 603 578 800 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=37640 $D=1
M708 606 569 604 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=33010 $D=1
M709 607 570 605 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=37640 $D=1
M710 604 577 606 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=33010 $D=1
M711 605 578 607 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=37640 $D=1
M712 6 602 604 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=33010 $D=1
M713 7 603 605 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=37640 $D=1
M714 608 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=33010 $D=1
M715 609 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=37640 $D=1
M716 610 608 596 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=33010 $D=1
M717 611 609 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=37640 $D=1
M718 600 129 610 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=33010 $D=1
M719 601 129 611 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=37640 $D=1
M720 612 608 598 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=33010 $D=1
M721 613 609 599 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=37640 $D=1
M722 606 129 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=33010 $D=1
M723 607 129 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=37640 $D=1
M724 614 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=33010 $D=1
M725 615 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=37640 $D=1
M726 616 614 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=33010 $D=1
M727 617 615 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=37640 $D=1
M728 610 130 616 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=33010 $D=1
M729 611 130 617 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=37640 $D=1
M730 14 616 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=33010 $D=1
M731 15 617 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=37640 $D=1
M732 618 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=33010 $D=1
M733 619 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=37640 $D=1
M734 620 618 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=33010 $D=1
M735 621 619 133 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=37640 $D=1
M736 134 131 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=33010 $D=1
M737 135 131 621 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=37640 $D=1
M738 622 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=33010 $D=1
M739 623 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=37640 $D=1
M740 624 622 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=33010 $D=1
M741 625 623 137 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=37640 $D=1
M742 138 131 624 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=33010 $D=1
M743 139 131 625 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=37640 $D=1
M744 626 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=33010 $D=1
M745 627 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=37640 $D=1
M746 628 626 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=33010 $D=1
M747 629 627 128 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=37640 $D=1
M748 140 131 628 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=33010 $D=1
M749 109 131 629 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=37640 $D=1
M750 630 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=33010 $D=1
M751 631 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=37640 $D=1
M752 632 630 141 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=33010 $D=1
M753 633 631 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=37640 $D=1
M754 143 131 632 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=33010 $D=1
M755 144 131 633 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=37640 $D=1
M756 634 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=33010 $D=1
M757 635 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=37640 $D=1
M758 636 634 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=33010 $D=1
M759 637 635 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=37640 $D=1
M760 143 131 636 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=33010 $D=1
M761 143 131 637 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=37640 $D=1
M762 6 569 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=33010 $D=1
M763 7 570 780 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=37640 $D=1
M764 135 779 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=33010 $D=1
M765 132 780 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=37640 $D=1
M766 638 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=33010 $D=1
M767 639 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=37640 $D=1
M768 148 638 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=33010 $D=1
M769 149 639 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=37640 $D=1
M770 620 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=33010 $D=1
M771 621 147 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=37640 $D=1
M772 640 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=33010 $D=1
M773 641 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=37640 $D=1
M774 151 640 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=33010 $D=1
M775 107 641 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=37640 $D=1
M776 624 150 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=33010 $D=1
M777 625 150 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=37640 $D=1
M778 642 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=33010 $D=1
M779 643 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=37640 $D=1
M780 153 642 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=33010 $D=1
M781 107 643 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=37640 $D=1
M782 628 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=33010 $D=1
M783 629 152 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=37640 $D=1
M784 644 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=33010 $D=1
M785 645 154 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=37640 $D=1
M786 155 644 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=33010 $D=1
M787 156 645 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=37640 $D=1
M788 632 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=33010 $D=1
M789 633 154 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=37640 $D=1
M790 646 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=33010 $D=1
M791 647 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=37640 $D=1
M792 219 646 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=33010 $D=1
M793 220 647 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=37640 $D=1
M794 636 157 219 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=33010 $D=1
M795 637 157 220 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=37640 $D=1
M796 648 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=33010 $D=1
M797 649 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=37640 $D=1
M798 650 648 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=33010 $D=1
M799 651 649 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=37640 $D=1
M800 12 158 650 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=33010 $D=1
M801 13 158 651 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=37640 $D=1
M802 801 559 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=33010 $D=1
M803 802 560 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=37640 $D=1
M804 652 650 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=33010 $D=1
M805 653 651 802 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=37640 $D=1
M806 656 559 654 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=33010 $D=1
M807 657 560 655 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=37640 $D=1
M808 654 650 656 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=33010 $D=1
M809 655 651 657 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=37640 $D=1
M810 6 652 654 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=33010 $D=1
M811 7 653 655 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=37640 $D=1
M812 803 159 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=33010 $D=1
M813 804 658 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=37640 $D=1
M814 781 656 803 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=33010 $D=1
M815 782 657 804 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=37640 $D=1
M816 658 781 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=33010 $D=1
M817 160 782 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=37640 $D=1
M818 659 559 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=33010 $D=1
M819 660 560 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=37640 $D=1
M820 6 661 659 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=33010 $D=1
M821 7 662 660 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=37640 $D=1
M822 661 650 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=33010 $D=1
M823 662 651 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=37640 $D=1
M824 805 659 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=33010 $D=1
M825 806 660 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=37640 $D=1
M826 663 159 805 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=33010 $D=1
M827 664 658 806 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=37640 $D=1
M828 666 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=33010 $D=1
M829 667 665 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=37640 $D=1
M830 807 663 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=33010 $D=1
M831 808 664 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=37640 $D=1
M832 665 666 807 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=33010 $D=1
M833 162 667 808 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=37640 $D=1
M834 669 668 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=33010 $D=1
M835 670 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=37640 $D=1
M836 6 673 671 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=33010 $D=1
M837 7 674 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=37640 $D=1
M838 675 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=33010 $D=1
M839 676 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=37640 $D=1
M840 673 675 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=33010 $D=1
M841 674 676 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=37640 $D=1
M842 669 121 673 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=33010 $D=1
M843 670 122 674 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=37640 $D=1
M844 677 671 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=33010 $D=1
M845 678 672 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=37640 $D=1
M846 164 677 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=33010 $D=1
M847 668 678 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=37640 $D=1
M848 121 671 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=33010 $D=1
M849 122 672 668 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=37640 $D=1
M850 679 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=33010 $D=1
M851 680 668 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=37640 $D=1
M852 681 671 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=33010 $D=1
M853 682 672 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=37640 $D=1
M854 221 681 679 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=33010 $D=1
M855 222 682 680 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=37640 $D=1
M856 6 671 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=33010 $D=1
M857 7 672 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=37640 $D=1
M858 683 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=33010 $D=1
M859 684 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=37640 $D=1
M860 685 683 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=33010 $D=1
M861 686 684 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=37640 $D=1
M862 14 165 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=33010 $D=1
M863 15 165 686 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=37640 $D=1
M864 687 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=33010 $D=1
M865 688 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=37640 $D=1
M866 166 687 685 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=33010 $D=1
M867 166 688 686 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=37640 $D=1
M868 6 166 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=33010 $D=1
M869 7 166 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=37640 $D=1
M870 689 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=33010 $D=1
M871 690 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=37640 $D=1
M872 6 689 691 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=33010 $D=1
M873 7 690 692 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=37640 $D=1
M874 693 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=33010 $D=1
M875 694 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=37640 $D=1
M876 695 689 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=33010 $D=1
M877 696 690 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=37640 $D=1
M878 6 695 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=33010 $D=1
M879 7 696 784 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=37640 $D=1
M880 697 783 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=33010 $D=1
M881 698 784 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=37640 $D=1
M882 695 691 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=33010 $D=1
M883 696 692 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=37640 $D=1
M884 699 117 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=33010 $D=1
M885 700 117 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=37640 $D=1
M886 6 703 701 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=33010 $D=1
M887 7 704 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=37640 $D=1
M888 703 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=33010 $D=1
M889 704 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=37640 $D=1
M890 785 699 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=33010 $D=1
M891 786 700 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=37640 $D=1
M892 705 701 785 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=33010 $D=1
M893 706 702 786 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=37640 $D=1
M894 6 705 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=33010 $D=1
M895 7 706 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=37640 $D=1
M896 787 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=33010 $D=1
M897 788 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=37640 $D=1
M898 705 703 787 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=33010 $D=1
M899 706 704 788 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=37640 $D=1
M900 195 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=34260 $D=0
M901 196 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=38890 $D=0
M902 197 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=34260 $D=0
M903 198 1 3 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=38890 $D=0
M904 6 195 197 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=34260 $D=0
M905 7 196 198 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=38890 $D=0
M906 199 1 4 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=34260 $D=0
M907 200 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=38890 $D=0
M908 5 195 199 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=34260 $D=0
M909 5 196 200 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=38890 $D=0
M910 201 1 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=34260 $D=0
M911 202 1 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=38890 $D=0
M912 6 195 201 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=34260 $D=0
M913 7 196 202 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=38890 $D=0
M914 205 9 201 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=34260 $D=0
M915 206 9 202 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=38890 $D=0
M916 203 9 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=34260 $D=0
M917 204 9 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=38890 $D=0
M918 207 9 199 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=34260 $D=0
M919 208 9 200 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=38890 $D=0
M920 197 203 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=34260 $D=0
M921 198 204 208 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=38890 $D=0
M922 209 10 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=34260 $D=0
M923 210 10 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=38890 $D=0
M924 211 10 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=34260 $D=0
M925 212 10 208 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=38890 $D=0
M926 205 209 211 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=34260 $D=0
M927 206 210 212 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=38890 $D=0
M928 213 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=34260 $D=0
M929 214 11 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=38890 $D=0
M930 215 11 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=34260 $D=0
M931 216 11 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=38890 $D=0
M932 12 213 215 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=34260 $D=0
M933 13 214 216 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=38890 $D=0
M934 217 11 14 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=34260 $D=0
M935 218 11 15 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=38890 $D=0
M936 219 213 217 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=34260 $D=0
M937 220 214 218 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=38890 $D=0
M938 223 11 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=34260 $D=0
M939 224 11 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=38890 $D=0
M940 211 213 223 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=34260 $D=0
M941 212 214 224 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=38890 $D=0
M942 227 16 223 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=34260 $D=0
M943 228 16 224 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=38890 $D=0
M944 225 16 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=34260 $D=0
M945 226 16 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=38890 $D=0
M946 229 16 217 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=34260 $D=0
M947 230 16 218 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=38890 $D=0
M948 215 225 229 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=34260 $D=0
M949 216 226 230 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=38890 $D=0
M950 231 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=34260 $D=0
M951 232 17 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=38890 $D=0
M952 233 17 229 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=34260 $D=0
M953 234 17 230 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=38890 $D=0
M954 227 231 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=34260 $D=0
M955 228 232 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=38890 $D=0
M956 167 18 235 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=34260 $D=0
M957 168 18 236 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=38890 $D=0
M958 237 19 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=34260 $D=0
M959 238 19 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=38890 $D=0
M960 239 235 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=34260 $D=0
M961 240 236 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=38890 $D=0
M962 167 239 707 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=34260 $D=0
M963 168 240 708 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=38890 $D=0
M964 241 707 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=34260 $D=0
M965 242 708 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=38890 $D=0
M966 239 18 241 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=34260 $D=0
M967 240 18 242 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=38890 $D=0
M968 241 237 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=34260 $D=0
M969 242 238 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=38890 $D=0
M970 247 245 241 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=34260 $D=0
M971 248 246 242 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=38890 $D=0
M972 245 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=34260 $D=0
M973 246 20 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=38890 $D=0
M974 167 21 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=34260 $D=0
M975 168 21 250 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=38890 $D=0
M976 251 22 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=34260 $D=0
M977 252 22 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=38890 $D=0
M978 253 249 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=34260 $D=0
M979 254 250 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=38890 $D=0
M980 167 253 709 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=34260 $D=0
M981 168 254 710 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=38890 $D=0
M982 255 709 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=34260 $D=0
M983 256 710 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=38890 $D=0
M984 253 21 255 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=34260 $D=0
M985 254 21 256 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=38890 $D=0
M986 255 251 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=34260 $D=0
M987 256 252 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=38890 $D=0
M988 247 257 255 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=34260 $D=0
M989 248 258 256 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=38890 $D=0
M990 257 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=34260 $D=0
M991 258 23 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=38890 $D=0
M992 167 24 259 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=34260 $D=0
M993 168 24 260 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=38890 $D=0
M994 261 25 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=34260 $D=0
M995 262 25 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=38890 $D=0
M996 263 259 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=34260 $D=0
M997 264 260 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=38890 $D=0
M998 167 263 711 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=34260 $D=0
M999 168 264 712 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=38890 $D=0
M1000 265 711 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=34260 $D=0
M1001 266 712 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=38890 $D=0
M1002 263 24 265 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=34260 $D=0
M1003 264 24 266 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=38890 $D=0
M1004 265 261 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=34260 $D=0
M1005 266 262 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=38890 $D=0
M1006 247 267 265 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=34260 $D=0
M1007 248 268 266 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=38890 $D=0
M1008 267 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=34260 $D=0
M1009 268 26 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=38890 $D=0
M1010 167 27 269 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=34260 $D=0
M1011 168 27 270 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=38890 $D=0
M1012 271 28 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=34260 $D=0
M1013 272 28 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=38890 $D=0
M1014 273 269 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=34260 $D=0
M1015 274 270 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=38890 $D=0
M1016 167 273 713 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=34260 $D=0
M1017 168 274 714 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=38890 $D=0
M1018 275 713 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=34260 $D=0
M1019 276 714 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=38890 $D=0
M1020 273 27 275 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=34260 $D=0
M1021 274 27 276 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=38890 $D=0
M1022 275 271 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=34260 $D=0
M1023 276 272 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=38890 $D=0
M1024 247 277 275 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=34260 $D=0
M1025 248 278 276 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=38890 $D=0
M1026 277 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=34260 $D=0
M1027 278 29 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=38890 $D=0
M1028 167 30 279 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=34260 $D=0
M1029 168 30 280 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=38890 $D=0
M1030 281 31 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=34260 $D=0
M1031 282 31 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=38890 $D=0
M1032 283 279 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=34260 $D=0
M1033 284 280 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=38890 $D=0
M1034 167 283 715 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=34260 $D=0
M1035 168 284 716 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=38890 $D=0
M1036 285 715 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=34260 $D=0
M1037 286 716 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=38890 $D=0
M1038 283 30 285 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=34260 $D=0
M1039 284 30 286 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=38890 $D=0
M1040 285 281 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=34260 $D=0
M1041 286 282 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=38890 $D=0
M1042 247 287 285 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=34260 $D=0
M1043 248 288 286 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=38890 $D=0
M1044 287 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=34260 $D=0
M1045 288 32 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=38890 $D=0
M1046 167 33 289 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=34260 $D=0
M1047 168 33 290 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=38890 $D=0
M1048 291 34 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=34260 $D=0
M1049 292 34 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=38890 $D=0
M1050 293 289 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=34260 $D=0
M1051 294 290 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=38890 $D=0
M1052 167 293 717 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=34260 $D=0
M1053 168 294 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=38890 $D=0
M1054 295 717 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=34260 $D=0
M1055 296 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=38890 $D=0
M1056 293 33 295 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=34260 $D=0
M1057 294 33 296 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=38890 $D=0
M1058 295 291 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=34260 $D=0
M1059 296 292 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=38890 $D=0
M1060 247 297 295 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=34260 $D=0
M1061 248 298 296 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=38890 $D=0
M1062 297 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=34260 $D=0
M1063 298 35 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=38890 $D=0
M1064 167 36 299 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=34260 $D=0
M1065 168 36 300 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=38890 $D=0
M1066 301 37 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=34260 $D=0
M1067 302 37 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=38890 $D=0
M1068 303 299 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=34260 $D=0
M1069 304 300 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=38890 $D=0
M1070 167 303 719 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=34260 $D=0
M1071 168 304 720 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=38890 $D=0
M1072 305 719 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=34260 $D=0
M1073 306 720 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=38890 $D=0
M1074 303 36 305 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=34260 $D=0
M1075 304 36 306 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=38890 $D=0
M1076 305 301 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=34260 $D=0
M1077 306 302 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=38890 $D=0
M1078 247 307 305 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=34260 $D=0
M1079 248 308 306 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=38890 $D=0
M1080 307 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=34260 $D=0
M1081 308 38 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=38890 $D=0
M1082 167 39 309 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=34260 $D=0
M1083 168 39 310 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=38890 $D=0
M1084 311 40 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=34260 $D=0
M1085 312 40 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=38890 $D=0
M1086 313 309 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=34260 $D=0
M1087 314 310 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=38890 $D=0
M1088 167 313 721 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=34260 $D=0
M1089 168 314 722 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=38890 $D=0
M1090 315 721 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=34260 $D=0
M1091 316 722 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=38890 $D=0
M1092 313 39 315 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=34260 $D=0
M1093 314 39 316 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=38890 $D=0
M1094 315 311 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=34260 $D=0
M1095 316 312 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=38890 $D=0
M1096 247 317 315 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=34260 $D=0
M1097 248 318 316 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=38890 $D=0
M1098 317 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=34260 $D=0
M1099 318 41 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=38890 $D=0
M1100 167 42 319 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=34260 $D=0
M1101 168 42 320 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=38890 $D=0
M1102 321 43 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=34260 $D=0
M1103 322 43 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=38890 $D=0
M1104 323 319 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=34260 $D=0
M1105 324 320 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=38890 $D=0
M1106 167 323 723 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=34260 $D=0
M1107 168 324 724 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=38890 $D=0
M1108 325 723 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=34260 $D=0
M1109 326 724 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=38890 $D=0
M1110 323 42 325 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=34260 $D=0
M1111 324 42 326 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=38890 $D=0
M1112 325 321 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=34260 $D=0
M1113 326 322 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=38890 $D=0
M1114 247 327 325 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=34260 $D=0
M1115 248 328 326 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=38890 $D=0
M1116 327 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=34260 $D=0
M1117 328 44 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=38890 $D=0
M1118 167 45 329 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=34260 $D=0
M1119 168 45 330 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=38890 $D=0
M1120 331 46 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=34260 $D=0
M1121 332 46 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=38890 $D=0
M1122 333 329 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=34260 $D=0
M1123 334 330 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=38890 $D=0
M1124 167 333 725 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=34260 $D=0
M1125 168 334 726 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=38890 $D=0
M1126 335 725 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=34260 $D=0
M1127 336 726 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=38890 $D=0
M1128 333 45 335 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=34260 $D=0
M1129 334 45 336 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=38890 $D=0
M1130 335 331 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=34260 $D=0
M1131 336 332 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=38890 $D=0
M1132 247 337 335 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=34260 $D=0
M1133 248 338 336 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=38890 $D=0
M1134 337 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=34260 $D=0
M1135 338 47 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=38890 $D=0
M1136 167 48 339 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=34260 $D=0
M1137 168 48 340 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=38890 $D=0
M1138 341 49 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=34260 $D=0
M1139 342 49 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=38890 $D=0
M1140 343 339 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=34260 $D=0
M1141 344 340 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=38890 $D=0
M1142 167 343 727 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=34260 $D=0
M1143 168 344 728 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=38890 $D=0
M1144 345 727 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=34260 $D=0
M1145 346 728 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=38890 $D=0
M1146 343 48 345 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=34260 $D=0
M1147 344 48 346 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=38890 $D=0
M1148 345 341 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=34260 $D=0
M1149 346 342 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=38890 $D=0
M1150 247 347 345 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=34260 $D=0
M1151 248 348 346 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=38890 $D=0
M1152 347 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=34260 $D=0
M1153 348 50 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=38890 $D=0
M1154 167 51 349 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=34260 $D=0
M1155 168 51 350 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=38890 $D=0
M1156 351 52 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=34260 $D=0
M1157 352 52 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=38890 $D=0
M1158 353 349 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=34260 $D=0
M1159 354 350 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=38890 $D=0
M1160 167 353 729 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=34260 $D=0
M1161 168 354 730 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=38890 $D=0
M1162 355 729 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=34260 $D=0
M1163 356 730 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=38890 $D=0
M1164 353 51 355 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=34260 $D=0
M1165 354 51 356 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=38890 $D=0
M1166 355 351 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=34260 $D=0
M1167 356 352 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=38890 $D=0
M1168 247 357 355 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=34260 $D=0
M1169 248 358 356 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=38890 $D=0
M1170 357 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=34260 $D=0
M1171 358 53 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=38890 $D=0
M1172 167 54 359 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=34260 $D=0
M1173 168 54 360 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=38890 $D=0
M1174 361 55 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=34260 $D=0
M1175 362 55 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=38890 $D=0
M1176 363 359 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=34260 $D=0
M1177 364 360 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=38890 $D=0
M1178 167 363 731 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=34260 $D=0
M1179 168 364 732 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=38890 $D=0
M1180 365 731 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=34260 $D=0
M1181 366 732 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=38890 $D=0
M1182 363 54 365 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=34260 $D=0
M1183 364 54 366 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=38890 $D=0
M1184 365 361 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=34260 $D=0
M1185 366 362 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=38890 $D=0
M1186 247 367 365 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=34260 $D=0
M1187 248 368 366 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=38890 $D=0
M1188 367 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=34260 $D=0
M1189 368 56 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=38890 $D=0
M1190 167 57 369 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=34260 $D=0
M1191 168 57 370 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=38890 $D=0
M1192 371 58 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=34260 $D=0
M1193 372 58 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=38890 $D=0
M1194 373 369 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=34260 $D=0
M1195 374 370 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=38890 $D=0
M1196 167 373 733 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=34260 $D=0
M1197 168 374 734 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=38890 $D=0
M1198 375 733 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=34260 $D=0
M1199 376 734 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=38890 $D=0
M1200 373 57 375 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=34260 $D=0
M1201 374 57 376 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=38890 $D=0
M1202 375 371 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=34260 $D=0
M1203 376 372 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=38890 $D=0
M1204 247 377 375 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=34260 $D=0
M1205 248 378 376 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=38890 $D=0
M1206 377 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=34260 $D=0
M1207 378 59 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=38890 $D=0
M1208 167 60 379 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=34260 $D=0
M1209 168 60 380 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=38890 $D=0
M1210 381 61 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=34260 $D=0
M1211 382 61 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=38890 $D=0
M1212 383 379 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=34260 $D=0
M1213 384 380 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=38890 $D=0
M1214 167 383 735 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=34260 $D=0
M1215 168 384 736 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=38890 $D=0
M1216 385 735 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=34260 $D=0
M1217 386 736 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=38890 $D=0
M1218 383 60 385 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=34260 $D=0
M1219 384 60 386 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=38890 $D=0
M1220 385 381 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=34260 $D=0
M1221 386 382 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=38890 $D=0
M1222 247 387 385 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=34260 $D=0
M1223 248 388 386 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=38890 $D=0
M1224 387 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=34260 $D=0
M1225 388 62 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=38890 $D=0
M1226 167 63 389 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=34260 $D=0
M1227 168 63 390 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=38890 $D=0
M1228 391 64 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=34260 $D=0
M1229 392 64 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=38890 $D=0
M1230 393 389 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=34260 $D=0
M1231 394 390 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=38890 $D=0
M1232 167 393 737 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=34260 $D=0
M1233 168 394 738 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=38890 $D=0
M1234 395 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=34260 $D=0
M1235 396 738 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=38890 $D=0
M1236 393 63 395 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=34260 $D=0
M1237 394 63 396 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=38890 $D=0
M1238 395 391 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=34260 $D=0
M1239 396 392 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=38890 $D=0
M1240 247 397 395 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=34260 $D=0
M1241 248 398 396 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=38890 $D=0
M1242 397 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=34260 $D=0
M1243 398 65 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=38890 $D=0
M1244 167 66 399 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=34260 $D=0
M1245 168 66 400 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=38890 $D=0
M1246 401 67 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=34260 $D=0
M1247 402 67 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=38890 $D=0
M1248 403 399 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=34260 $D=0
M1249 404 400 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=38890 $D=0
M1250 167 403 739 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=34260 $D=0
M1251 168 404 740 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=38890 $D=0
M1252 405 739 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=34260 $D=0
M1253 406 740 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=38890 $D=0
M1254 403 66 405 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=34260 $D=0
M1255 404 66 406 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=38890 $D=0
M1256 405 401 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=34260 $D=0
M1257 406 402 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=38890 $D=0
M1258 247 407 405 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=34260 $D=0
M1259 248 408 406 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=38890 $D=0
M1260 407 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=34260 $D=0
M1261 408 68 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=38890 $D=0
M1262 167 69 409 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=34260 $D=0
M1263 168 69 410 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=38890 $D=0
M1264 411 70 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=34260 $D=0
M1265 412 70 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=38890 $D=0
M1266 413 409 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=34260 $D=0
M1267 414 410 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=38890 $D=0
M1268 167 413 741 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=34260 $D=0
M1269 168 414 742 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=38890 $D=0
M1270 415 741 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=34260 $D=0
M1271 416 742 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=38890 $D=0
M1272 413 69 415 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=34260 $D=0
M1273 414 69 416 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=38890 $D=0
M1274 415 411 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=34260 $D=0
M1275 416 412 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=38890 $D=0
M1276 247 417 415 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=34260 $D=0
M1277 248 418 416 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=38890 $D=0
M1278 417 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=34260 $D=0
M1279 418 71 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=38890 $D=0
M1280 167 72 419 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=34260 $D=0
M1281 168 72 420 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=38890 $D=0
M1282 421 73 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=34260 $D=0
M1283 422 73 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=38890 $D=0
M1284 423 419 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=34260 $D=0
M1285 424 420 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=38890 $D=0
M1286 167 423 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=34260 $D=0
M1287 168 424 744 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=38890 $D=0
M1288 425 743 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=34260 $D=0
M1289 426 744 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=38890 $D=0
M1290 423 72 425 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=34260 $D=0
M1291 424 72 426 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=38890 $D=0
M1292 425 421 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=34260 $D=0
M1293 426 422 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=38890 $D=0
M1294 247 427 425 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=34260 $D=0
M1295 248 428 426 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=38890 $D=0
M1296 427 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=34260 $D=0
M1297 428 74 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=38890 $D=0
M1298 167 75 429 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=34260 $D=0
M1299 168 75 430 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=38890 $D=0
M1300 431 76 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=34260 $D=0
M1301 432 76 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=38890 $D=0
M1302 433 429 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=34260 $D=0
M1303 434 430 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=38890 $D=0
M1304 167 433 745 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=34260 $D=0
M1305 168 434 746 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=38890 $D=0
M1306 435 745 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=34260 $D=0
M1307 436 746 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=38890 $D=0
M1308 433 75 435 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=34260 $D=0
M1309 434 75 436 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=38890 $D=0
M1310 435 431 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=34260 $D=0
M1311 436 432 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=38890 $D=0
M1312 247 437 435 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=34260 $D=0
M1313 248 438 436 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=38890 $D=0
M1314 437 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=34260 $D=0
M1315 438 77 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=38890 $D=0
M1316 167 78 439 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=34260 $D=0
M1317 168 78 440 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=38890 $D=0
M1318 441 79 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=34260 $D=0
M1319 442 79 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=38890 $D=0
M1320 443 439 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=34260 $D=0
M1321 444 440 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=38890 $D=0
M1322 167 443 747 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=34260 $D=0
M1323 168 444 748 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=38890 $D=0
M1324 445 747 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=34260 $D=0
M1325 446 748 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=38890 $D=0
M1326 443 78 445 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=34260 $D=0
M1327 444 78 446 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=38890 $D=0
M1328 445 441 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=34260 $D=0
M1329 446 442 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=38890 $D=0
M1330 247 447 445 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=34260 $D=0
M1331 248 448 446 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=38890 $D=0
M1332 447 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=34260 $D=0
M1333 448 80 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=38890 $D=0
M1334 167 81 449 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=34260 $D=0
M1335 168 81 450 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=38890 $D=0
M1336 451 82 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=34260 $D=0
M1337 452 82 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=38890 $D=0
M1338 453 449 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=34260 $D=0
M1339 454 450 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=38890 $D=0
M1340 167 453 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=34260 $D=0
M1341 168 454 750 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=38890 $D=0
M1342 455 749 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=34260 $D=0
M1343 456 750 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=38890 $D=0
M1344 453 81 455 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=34260 $D=0
M1345 454 81 456 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=38890 $D=0
M1346 455 451 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=34260 $D=0
M1347 456 452 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=38890 $D=0
M1348 247 457 455 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=34260 $D=0
M1349 248 458 456 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=38890 $D=0
M1350 457 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=34260 $D=0
M1351 458 83 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=38890 $D=0
M1352 167 84 459 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=34260 $D=0
M1353 168 84 460 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=38890 $D=0
M1354 461 85 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=34260 $D=0
M1355 462 85 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=38890 $D=0
M1356 463 459 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=34260 $D=0
M1357 464 460 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=38890 $D=0
M1358 167 463 751 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=34260 $D=0
M1359 168 464 752 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=38890 $D=0
M1360 465 751 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=34260 $D=0
M1361 466 752 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=38890 $D=0
M1362 463 84 465 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=34260 $D=0
M1363 464 84 466 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=38890 $D=0
M1364 465 461 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=34260 $D=0
M1365 466 462 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=38890 $D=0
M1366 247 467 465 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=34260 $D=0
M1367 248 468 466 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=38890 $D=0
M1368 467 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=34260 $D=0
M1369 468 86 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=38890 $D=0
M1370 167 87 469 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=34260 $D=0
M1371 168 87 470 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=38890 $D=0
M1372 471 88 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=34260 $D=0
M1373 472 88 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=38890 $D=0
M1374 473 469 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=34260 $D=0
M1375 474 470 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=38890 $D=0
M1376 167 473 753 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=34260 $D=0
M1377 168 474 754 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=38890 $D=0
M1378 475 753 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=34260 $D=0
M1379 476 754 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=38890 $D=0
M1380 473 87 475 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=34260 $D=0
M1381 474 87 476 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=38890 $D=0
M1382 475 471 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=34260 $D=0
M1383 476 472 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=38890 $D=0
M1384 247 477 475 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=34260 $D=0
M1385 248 478 476 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=38890 $D=0
M1386 477 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=34260 $D=0
M1387 478 89 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=38890 $D=0
M1388 167 90 479 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=34260 $D=0
M1389 168 90 480 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=38890 $D=0
M1390 481 91 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=34260 $D=0
M1391 482 91 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=38890 $D=0
M1392 483 479 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=34260 $D=0
M1393 484 480 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=38890 $D=0
M1394 167 483 755 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=34260 $D=0
M1395 168 484 756 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=38890 $D=0
M1396 485 755 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=34260 $D=0
M1397 486 756 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=38890 $D=0
M1398 483 90 485 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=34260 $D=0
M1399 484 90 486 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=38890 $D=0
M1400 485 481 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=34260 $D=0
M1401 486 482 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=38890 $D=0
M1402 247 487 485 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=34260 $D=0
M1403 248 488 486 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=38890 $D=0
M1404 487 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=34260 $D=0
M1405 488 92 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=38890 $D=0
M1406 167 93 489 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=34260 $D=0
M1407 168 93 490 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=38890 $D=0
M1408 491 94 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=34260 $D=0
M1409 492 94 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=38890 $D=0
M1410 493 489 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=34260 $D=0
M1411 494 490 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=38890 $D=0
M1412 167 493 757 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=34260 $D=0
M1413 168 494 758 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=38890 $D=0
M1414 495 757 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=34260 $D=0
M1415 496 758 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=38890 $D=0
M1416 493 93 495 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=34260 $D=0
M1417 494 93 496 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=38890 $D=0
M1418 495 491 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=34260 $D=0
M1419 496 492 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=38890 $D=0
M1420 247 497 495 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=34260 $D=0
M1421 248 498 496 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=38890 $D=0
M1422 497 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=34260 $D=0
M1423 498 95 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=38890 $D=0
M1424 167 96 499 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=34260 $D=0
M1425 168 96 500 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=38890 $D=0
M1426 501 97 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=34260 $D=0
M1427 502 97 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=38890 $D=0
M1428 503 499 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=34260 $D=0
M1429 504 500 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=38890 $D=0
M1430 167 503 759 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=34260 $D=0
M1431 168 504 760 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=38890 $D=0
M1432 505 759 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=34260 $D=0
M1433 506 760 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=38890 $D=0
M1434 503 96 505 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=34260 $D=0
M1435 504 96 506 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=38890 $D=0
M1436 505 501 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=34260 $D=0
M1437 506 502 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=38890 $D=0
M1438 247 507 505 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=34260 $D=0
M1439 248 508 506 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=38890 $D=0
M1440 507 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=34260 $D=0
M1441 508 98 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=38890 $D=0
M1442 167 99 509 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=34260 $D=0
M1443 168 99 510 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=38890 $D=0
M1444 511 100 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=34260 $D=0
M1445 512 100 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=38890 $D=0
M1446 513 509 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=34260 $D=0
M1447 514 510 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=38890 $D=0
M1448 167 513 761 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=34260 $D=0
M1449 168 514 762 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=38890 $D=0
M1450 515 761 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=34260 $D=0
M1451 516 762 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=38890 $D=0
M1452 513 99 515 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=34260 $D=0
M1453 514 99 516 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=38890 $D=0
M1454 515 511 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=34260 $D=0
M1455 516 512 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=38890 $D=0
M1456 247 517 515 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=34260 $D=0
M1457 248 518 516 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=38890 $D=0
M1458 517 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=34260 $D=0
M1459 518 101 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=38890 $D=0
M1460 167 102 519 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=34260 $D=0
M1461 168 102 520 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=38890 $D=0
M1462 521 103 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=34260 $D=0
M1463 522 103 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=38890 $D=0
M1464 523 519 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=34260 $D=0
M1465 524 520 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=38890 $D=0
M1466 167 523 763 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=34260 $D=0
M1467 168 524 764 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=38890 $D=0
M1468 525 763 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=34260 $D=0
M1469 526 764 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=38890 $D=0
M1470 523 102 525 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=34260 $D=0
M1471 524 102 526 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=38890 $D=0
M1472 525 521 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=34260 $D=0
M1473 526 522 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=38890 $D=0
M1474 247 527 525 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=34260 $D=0
M1475 248 528 526 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=38890 $D=0
M1476 527 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=34260 $D=0
M1477 528 104 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=38890 $D=0
M1478 167 105 529 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=34260 $D=0
M1479 168 105 530 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=38890 $D=0
M1480 531 106 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=34260 $D=0
M1481 532 106 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=38890 $D=0
M1482 533 529 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=34260 $D=0
M1483 534 530 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=38890 $D=0
M1484 167 533 765 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=34260 $D=0
M1485 168 534 766 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=38890 $D=0
M1486 535 765 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=34260 $D=0
M1487 536 766 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=38890 $D=0
M1488 533 105 535 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=34260 $D=0
M1489 534 105 536 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=38890 $D=0
M1490 535 531 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=34260 $D=0
M1491 536 532 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=38890 $D=0
M1492 247 537 535 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=34260 $D=0
M1493 248 538 536 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=38890 $D=0
M1494 537 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=34260 $D=0
M1495 538 110 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=38890 $D=0
M1496 167 112 539 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=34260 $D=0
M1497 168 112 540 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=38890 $D=0
M1498 541 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=34260 $D=0
M1499 542 113 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=38890 $D=0
M1500 543 539 233 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=34260 $D=0
M1501 544 540 234 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=38890 $D=0
M1502 167 543 767 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=34260 $D=0
M1503 168 544 768 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=38890 $D=0
M1504 545 767 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=34260 $D=0
M1505 546 768 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=38890 $D=0
M1506 543 112 545 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=34260 $D=0
M1507 544 112 546 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=38890 $D=0
M1508 545 541 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=34260 $D=0
M1509 546 542 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=38890 $D=0
M1510 247 547 545 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=34260 $D=0
M1511 248 548 546 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=38890 $D=0
M1512 547 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=34260 $D=0
M1513 548 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=38890 $D=0
M1514 167 115 549 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=34260 $D=0
M1515 168 115 550 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=38890 $D=0
M1516 551 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=34260 $D=0
M1517 552 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=38890 $D=0
M1518 6 551 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=34260 $D=0
M1519 7 552 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=38890 $D=0
M1520 247 549 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=34260 $D=0
M1521 248 550 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=38890 $D=0
M1522 167 555 553 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=34260 $D=0
M1523 168 556 554 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=38890 $D=0
M1524 555 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=34260 $D=0
M1525 556 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=38890 $D=0
M1526 769 243 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=34260 $D=0
M1527 770 244 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=38890 $D=0
M1528 557 555 769 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=34260 $D=0
M1529 558 556 770 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=38890 $D=0
M1530 167 557 559 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=34260 $D=0
M1531 168 558 560 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=38890 $D=0
M1532 771 559 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=34260 $D=0
M1533 772 560 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=38890 $D=0
M1534 557 553 771 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=34260 $D=0
M1535 558 554 772 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=38890 $D=0
M1536 167 563 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=34260 $D=0
M1537 168 564 562 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=38890 $D=0
M1538 563 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=34260 $D=0
M1539 564 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=38890 $D=0
M1540 773 247 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=34260 $D=0
M1541 774 248 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=38890 $D=0
M1542 565 563 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=34260 $D=0
M1543 566 564 774 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=38890 $D=0
M1544 167 565 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=34260 $D=0
M1545 168 566 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=38890 $D=0
M1546 775 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=34260 $D=0
M1547 776 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=38890 $D=0
M1548 565 561 775 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=34260 $D=0
M1549 566 562 776 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=38890 $D=0
M1550 567 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=34260 $D=0
M1551 568 120 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=38890 $D=0
M1552 569 120 559 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=34260 $D=0
M1553 570 120 560 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=38890 $D=0
M1554 121 567 569 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=34260 $D=0
M1555 122 568 570 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=38890 $D=0
M1556 571 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=34260 $D=0
M1557 572 123 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=38890 $D=0
M1558 573 123 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=34260 $D=0
M1559 574 123 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=38890 $D=0
M1560 777 571 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=34260 $D=0
M1561 778 572 574 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=38890 $D=0
M1562 167 118 777 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=34260 $D=0
M1563 168 119 778 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=38890 $D=0
M1564 575 124 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=34260 $D=0
M1565 576 124 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=38890 $D=0
M1566 577 124 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=34260 $D=0
M1567 578 124 574 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=38890 $D=0
M1568 12 575 577 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=34260 $D=0
M1569 13 576 578 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=38890 $D=0
M1570 580 579 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=34260 $D=0
M1571 581 125 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=38890 $D=0
M1572 167 584 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=34260 $D=0
M1573 168 585 583 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=38890 $D=0
M1574 586 569 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=34260 $D=0
M1575 587 570 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=38890 $D=0
M1576 584 569 579 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=34260 $D=0
M1577 585 570 125 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=38890 $D=0
M1578 580 586 584 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=34260 $D=0
M1579 581 587 585 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=38890 $D=0
M1580 588 582 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=34260 $D=0
M1581 589 583 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=38890 $D=0
M1582 126 582 577 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=34260 $D=0
M1583 579 583 578 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=38890 $D=0
M1584 569 588 126 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=34260 $D=0
M1585 570 589 579 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=38890 $D=0
M1586 590 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=34260 $D=0
M1587 591 579 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=38890 $D=0
M1588 592 582 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=34260 $D=0
M1589 593 583 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=38890 $D=0
M1590 594 582 590 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=34260 $D=0
M1591 595 583 591 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=38890 $D=0
M1592 577 592 594 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=34260 $D=0
M1593 578 593 595 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=38890 $D=0
M1594 789 569 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=33900 $D=0
M1595 790 570 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=38530 $D=0
M1596 596 577 789 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=33900 $D=0
M1597 597 578 790 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=38530 $D=0
M1598 598 594 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=34260 $D=0
M1599 599 595 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=38890 $D=0
M1600 600 569 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=34260 $D=0
M1601 601 570 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=38890 $D=0
M1602 167 577 600 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=34260 $D=0
M1603 168 578 601 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=38890 $D=0
M1604 602 569 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=34260 $D=0
M1605 603 570 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=38890 $D=0
M1606 167 577 602 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=34260 $D=0
M1607 168 578 603 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=38890 $D=0
M1608 791 569 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=34080 $D=0
M1609 792 570 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=38710 $D=0
M1610 606 577 791 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=34080 $D=0
M1611 607 578 792 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=38710 $D=0
M1612 167 602 606 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=34260 $D=0
M1613 168 603 607 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=38890 $D=0
M1614 608 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=34260 $D=0
M1615 609 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=38890 $D=0
M1616 610 129 596 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=34260 $D=0
M1617 611 129 597 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=38890 $D=0
M1618 600 608 610 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=34260 $D=0
M1619 601 609 611 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=38890 $D=0
M1620 612 129 598 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=34260 $D=0
M1621 613 129 599 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=38890 $D=0
M1622 606 608 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=34260 $D=0
M1623 607 609 613 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=38890 $D=0
M1624 614 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=34260 $D=0
M1625 615 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=38890 $D=0
M1626 616 130 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=34260 $D=0
M1627 617 130 613 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=38890 $D=0
M1628 610 614 616 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=34260 $D=0
M1629 611 615 617 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=38890 $D=0
M1630 14 616 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=34260 $D=0
M1631 15 617 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=38890 $D=0
M1632 618 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=34260 $D=0
M1633 619 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=38890 $D=0
M1634 620 131 132 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=34260 $D=0
M1635 621 131 133 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=38890 $D=0
M1636 134 618 620 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=34260 $D=0
M1637 135 619 621 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=38890 $D=0
M1638 622 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=34260 $D=0
M1639 623 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=38890 $D=0
M1640 624 131 136 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=34260 $D=0
M1641 625 131 137 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=38890 $D=0
M1642 138 622 624 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=34260 $D=0
M1643 139 623 625 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=38890 $D=0
M1644 626 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=34260 $D=0
M1645 627 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=38890 $D=0
M1646 628 131 127 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=34260 $D=0
M1647 629 131 128 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=38890 $D=0
M1648 140 626 628 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=34260 $D=0
M1649 109 627 629 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=38890 $D=0
M1650 630 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=34260 $D=0
M1651 631 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=38890 $D=0
M1652 632 131 141 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=34260 $D=0
M1653 633 131 142 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=38890 $D=0
M1654 143 630 632 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=34260 $D=0
M1655 144 631 633 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=38890 $D=0
M1656 634 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=34260 $D=0
M1657 635 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=38890 $D=0
M1658 636 131 145 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=34260 $D=0
M1659 637 131 146 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=38890 $D=0
M1660 143 634 636 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=34260 $D=0
M1661 143 635 637 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=38890 $D=0
M1662 167 569 779 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=34260 $D=0
M1663 168 570 780 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=38890 $D=0
M1664 135 779 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=34260 $D=0
M1665 132 780 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=38890 $D=0
M1666 638 147 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=34260 $D=0
M1667 639 147 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=38890 $D=0
M1668 148 147 135 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=34260 $D=0
M1669 149 147 132 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=38890 $D=0
M1670 620 638 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=34260 $D=0
M1671 621 639 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=38890 $D=0
M1672 640 150 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=34260 $D=0
M1673 641 150 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=38890 $D=0
M1674 151 150 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=34260 $D=0
M1675 107 150 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=38890 $D=0
M1676 624 640 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=34260 $D=0
M1677 625 641 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=38890 $D=0
M1678 642 152 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=34260 $D=0
M1679 643 152 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=38890 $D=0
M1680 153 152 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=34260 $D=0
M1681 107 152 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=38890 $D=0
M1682 628 642 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=34260 $D=0
M1683 629 643 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=38890 $D=0
M1684 644 154 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=34260 $D=0
M1685 645 154 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=38890 $D=0
M1686 155 154 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=34260 $D=0
M1687 156 154 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=38890 $D=0
M1688 632 644 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=34260 $D=0
M1689 633 645 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=38890 $D=0
M1690 646 157 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=34260 $D=0
M1691 647 157 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=38890 $D=0
M1692 219 157 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=34260 $D=0
M1693 220 157 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=38890 $D=0
M1694 636 646 219 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=34260 $D=0
M1695 637 647 220 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=38890 $D=0
M1696 648 158 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=34260 $D=0
M1697 649 158 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=38890 $D=0
M1698 650 158 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=34260 $D=0
M1699 651 158 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=38890 $D=0
M1700 12 648 650 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=34260 $D=0
M1701 13 649 651 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=38890 $D=0
M1702 652 559 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=34260 $D=0
M1703 653 560 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=38890 $D=0
M1704 167 650 652 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=34260 $D=0
M1705 168 651 653 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=38890 $D=0
M1706 793 559 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=34080 $D=0
M1707 794 560 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=38710 $D=0
M1708 656 650 793 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=34080 $D=0
M1709 657 651 794 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=38710 $D=0
M1710 167 652 656 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=34260 $D=0
M1711 168 653 657 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=38890 $D=0
M1712 781 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=34260 $D=0
M1713 782 658 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=38890 $D=0
M1714 167 656 781 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=34260 $D=0
M1715 168 657 782 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=38890 $D=0
M1716 658 781 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=34260 $D=0
M1717 160 782 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=38890 $D=0
M1718 795 559 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=33900 $D=0
M1719 796 560 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=38530 $D=0
M1720 659 661 795 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=33900 $D=0
M1721 660 662 796 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=38530 $D=0
M1722 661 650 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=34260 $D=0
M1723 662 651 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=38890 $D=0
M1724 663 659 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=34260 $D=0
M1725 664 660 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=38890 $D=0
M1726 167 159 663 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=34260 $D=0
M1727 168 658 664 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=38890 $D=0
M1728 666 161 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=34260 $D=0
M1729 667 665 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=38890 $D=0
M1730 665 663 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=34260 $D=0
M1731 162 664 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=38890 $D=0
M1732 167 666 665 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=34260 $D=0
M1733 168 667 162 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=38890 $D=0
M1734 669 668 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=34260 $D=0
M1735 670 163 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=38890 $D=0
M1736 167 673 671 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=34260 $D=0
M1737 168 674 672 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=38890 $D=0
M1738 675 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=34260 $D=0
M1739 676 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=38890 $D=0
M1740 673 121 668 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=34260 $D=0
M1741 674 122 163 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=38890 $D=0
M1742 669 675 673 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=34260 $D=0
M1743 670 676 674 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=38890 $D=0
M1744 677 671 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=34260 $D=0
M1745 678 672 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=38890 $D=0
M1746 164 671 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=34260 $D=0
M1747 668 672 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=38890 $D=0
M1748 121 677 164 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=34260 $D=0
M1749 122 678 668 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=38890 $D=0
M1750 679 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=34260 $D=0
M1751 680 668 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=38890 $D=0
M1752 681 671 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=34260 $D=0
M1753 682 672 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=38890 $D=0
M1754 221 671 679 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=34260 $D=0
M1755 222 672 680 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=38890 $D=0
M1756 6 681 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=34260 $D=0
M1757 7 682 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=38890 $D=0
M1758 683 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=34260 $D=0
M1759 684 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=38890 $D=0
M1760 685 165 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=34260 $D=0
M1761 686 165 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=38890 $D=0
M1762 14 683 685 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=34260 $D=0
M1763 15 684 686 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=38890 $D=0
M1764 687 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=34260 $D=0
M1765 688 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=38890 $D=0
M1766 166 166 685 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=34260 $D=0
M1767 166 166 686 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=38890 $D=0
M1768 6 687 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=34260 $D=0
M1769 7 688 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=38890 $D=0
M1770 689 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=34260 $D=0
M1771 690 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=38890 $D=0
M1772 167 689 691 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=34260 $D=0
M1773 168 690 692 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=38890 $D=0
M1774 693 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=34260 $D=0
M1775 694 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=38890 $D=0
M1776 695 691 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=34260 $D=0
M1777 696 692 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=38890 $D=0
M1778 167 695 783 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=34260 $D=0
M1779 168 696 784 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=38890 $D=0
M1780 697 783 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=34260 $D=0
M1781 698 784 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=38890 $D=0
M1782 695 689 697 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=34260 $D=0
M1783 696 690 698 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=38890 $D=0
M1784 699 693 697 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=34260 $D=0
M1785 700 694 698 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=38890 $D=0
M1786 167 703 701 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=34260 $D=0
M1787 168 704 702 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=38890 $D=0
M1788 703 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=34260 $D=0
M1789 704 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=38890 $D=0
M1790 785 699 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=34260 $D=0
M1791 786 700 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=38890 $D=0
M1792 705 703 785 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=34260 $D=0
M1793 706 704 786 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=38890 $D=0
M1794 167 705 121 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=34260 $D=0
M1795 168 706 122 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=38890 $D=0
M1796 787 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=34260 $D=0
M1797 788 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=38890 $D=0
M1798 705 701 787 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=34260 $D=0
M1799 706 702 788 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=38890 $D=0
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 112 113 114 115 116 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168
** N=804 EP=164 IP=1514 FDC=1800
M0 190 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=23750 $D=1
M1 191 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=28380 $D=1
M2 192 190 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=23750 $D=1
M3 193 191 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=28380 $D=1
M4 6 1 192 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=23750 $D=1
M5 7 1 193 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=28380 $D=1
M6 194 190 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=23750 $D=1
M7 195 191 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=28380 $D=1
M8 5 1 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=23750 $D=1
M9 5 1 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=28380 $D=1
M10 196 190 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=23750 $D=1
M11 197 191 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=28380 $D=1
M12 6 1 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=23750 $D=1
M13 7 1 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=28380 $D=1
M14 200 198 196 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=23750 $D=1
M15 201 199 197 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=28380 $D=1
M16 198 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=23750 $D=1
M17 199 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=28380 $D=1
M18 202 198 194 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=23750 $D=1
M19 203 199 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=28380 $D=1
M20 192 9 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=23750 $D=1
M21 193 9 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=28380 $D=1
M22 204 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=23750 $D=1
M23 205 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=28380 $D=1
M24 206 204 202 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=23750 $D=1
M25 207 205 203 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=28380 $D=1
M26 200 10 206 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=23750 $D=1
M27 201 10 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=28380 $D=1
M28 208 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=23750 $D=1
M29 209 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=28380 $D=1
M30 210 208 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=23750 $D=1
M31 211 209 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=28380 $D=1
M32 12 11 210 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=23750 $D=1
M33 13 11 211 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=28380 $D=1
M34 212 208 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=23750 $D=1
M35 213 209 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=28380 $D=1
M36 214 11 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=23750 $D=1
M37 215 11 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=28380 $D=1
M38 218 208 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=23750 $D=1
M39 219 209 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=28380 $D=1
M40 206 11 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=23750 $D=1
M41 207 11 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=28380 $D=1
M42 222 220 218 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=23750 $D=1
M43 223 221 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=28380 $D=1
M44 220 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=23750 $D=1
M45 221 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=28380 $D=1
M46 224 220 212 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=23750 $D=1
M47 225 221 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=28380 $D=1
M48 210 16 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=23750 $D=1
M49 211 16 225 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=28380 $D=1
M50 226 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=23750 $D=1
M51 227 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=28380 $D=1
M52 228 226 224 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=23750 $D=1
M53 229 227 225 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=28380 $D=1
M54 222 17 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=23750 $D=1
M55 223 17 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=28380 $D=1
M56 6 18 230 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=23750 $D=1
M57 7 18 231 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=28380 $D=1
M58 232 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=23750 $D=1
M59 233 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=28380 $D=1
M60 234 18 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=23750 $D=1
M61 235 18 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=28380 $D=1
M62 6 234 703 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=23750 $D=1
M63 7 235 704 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=28380 $D=1
M64 236 703 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=23750 $D=1
M65 237 704 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=28380 $D=1
M66 234 230 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=23750 $D=1
M67 235 231 237 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=28380 $D=1
M68 236 19 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=23750 $D=1
M69 237 19 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=28380 $D=1
M70 242 20 236 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=23750 $D=1
M71 243 20 237 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=28380 $D=1
M72 240 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=23750 $D=1
M73 241 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=28380 $D=1
M74 6 21 244 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=23750 $D=1
M75 7 21 245 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=28380 $D=1
M76 246 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=23750 $D=1
M77 247 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=28380 $D=1
M78 248 21 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=23750 $D=1
M79 249 21 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=28380 $D=1
M80 6 248 705 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=23750 $D=1
M81 7 249 706 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=28380 $D=1
M82 250 705 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=23750 $D=1
M83 251 706 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=28380 $D=1
M84 248 244 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=23750 $D=1
M85 249 245 251 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=28380 $D=1
M86 250 22 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=23750 $D=1
M87 251 22 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=28380 $D=1
M88 242 23 250 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=23750 $D=1
M89 243 23 251 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=28380 $D=1
M90 252 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=23750 $D=1
M91 253 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=28380 $D=1
M92 6 24 254 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=23750 $D=1
M93 7 24 255 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=28380 $D=1
M94 256 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=23750 $D=1
M95 257 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=28380 $D=1
M96 258 24 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=23750 $D=1
M97 259 24 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=28380 $D=1
M98 6 258 707 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=23750 $D=1
M99 7 259 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=28380 $D=1
M100 260 707 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=23750 $D=1
M101 261 708 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=28380 $D=1
M102 258 254 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=23750 $D=1
M103 259 255 261 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=28380 $D=1
M104 260 25 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=23750 $D=1
M105 261 25 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=28380 $D=1
M106 242 26 260 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=23750 $D=1
M107 243 26 261 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=28380 $D=1
M108 262 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=23750 $D=1
M109 263 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=28380 $D=1
M110 6 27 264 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=23750 $D=1
M111 7 27 265 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=28380 $D=1
M112 266 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=23750 $D=1
M113 267 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=28380 $D=1
M114 268 27 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=23750 $D=1
M115 269 27 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=28380 $D=1
M116 6 268 709 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=23750 $D=1
M117 7 269 710 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=28380 $D=1
M118 270 709 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=23750 $D=1
M119 271 710 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=28380 $D=1
M120 268 264 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=23750 $D=1
M121 269 265 271 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=28380 $D=1
M122 270 28 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=23750 $D=1
M123 271 28 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=28380 $D=1
M124 242 29 270 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=23750 $D=1
M125 243 29 271 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=28380 $D=1
M126 272 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=23750 $D=1
M127 273 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=28380 $D=1
M128 6 30 274 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=23750 $D=1
M129 7 30 275 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=28380 $D=1
M130 276 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=23750 $D=1
M131 277 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=28380 $D=1
M132 278 30 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=23750 $D=1
M133 279 30 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=28380 $D=1
M134 6 278 711 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=23750 $D=1
M135 7 279 712 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=28380 $D=1
M136 280 711 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=23750 $D=1
M137 281 712 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=28380 $D=1
M138 278 274 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=23750 $D=1
M139 279 275 281 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=28380 $D=1
M140 280 31 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=23750 $D=1
M141 281 31 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=28380 $D=1
M142 242 32 280 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=23750 $D=1
M143 243 32 281 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=28380 $D=1
M144 282 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=23750 $D=1
M145 283 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=28380 $D=1
M146 6 33 284 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=23750 $D=1
M147 7 33 285 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=28380 $D=1
M148 286 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=23750 $D=1
M149 287 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=28380 $D=1
M150 288 33 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=23750 $D=1
M151 289 33 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=28380 $D=1
M152 6 288 713 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=23750 $D=1
M153 7 289 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=28380 $D=1
M154 290 713 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=23750 $D=1
M155 291 714 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=28380 $D=1
M156 288 284 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=23750 $D=1
M157 289 285 291 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=28380 $D=1
M158 290 34 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=23750 $D=1
M159 291 34 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=28380 $D=1
M160 242 35 290 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=23750 $D=1
M161 243 35 291 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=28380 $D=1
M162 292 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=23750 $D=1
M163 293 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=28380 $D=1
M164 6 36 294 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=23750 $D=1
M165 7 36 295 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=28380 $D=1
M166 296 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=23750 $D=1
M167 297 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=28380 $D=1
M168 298 36 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=23750 $D=1
M169 299 36 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=28380 $D=1
M170 6 298 715 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=23750 $D=1
M171 7 299 716 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=28380 $D=1
M172 300 715 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=23750 $D=1
M173 301 716 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=28380 $D=1
M174 298 294 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=23750 $D=1
M175 299 295 301 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=28380 $D=1
M176 300 37 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=23750 $D=1
M177 301 37 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=28380 $D=1
M178 242 38 300 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=23750 $D=1
M179 243 38 301 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=28380 $D=1
M180 302 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=23750 $D=1
M181 303 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=28380 $D=1
M182 6 39 304 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=23750 $D=1
M183 7 39 305 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=28380 $D=1
M184 306 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=23750 $D=1
M185 307 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=28380 $D=1
M186 308 39 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=23750 $D=1
M187 309 39 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=28380 $D=1
M188 6 308 717 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=23750 $D=1
M189 7 309 718 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=28380 $D=1
M190 310 717 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=23750 $D=1
M191 311 718 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=28380 $D=1
M192 308 304 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=23750 $D=1
M193 309 305 311 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=28380 $D=1
M194 310 40 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=23750 $D=1
M195 311 40 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=28380 $D=1
M196 242 41 310 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=23750 $D=1
M197 243 41 311 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=28380 $D=1
M198 312 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=23750 $D=1
M199 313 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=28380 $D=1
M200 6 42 314 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=23750 $D=1
M201 7 42 315 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=28380 $D=1
M202 316 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=23750 $D=1
M203 317 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=28380 $D=1
M204 318 42 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=23750 $D=1
M205 319 42 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=28380 $D=1
M206 6 318 719 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=23750 $D=1
M207 7 319 720 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=28380 $D=1
M208 320 719 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=23750 $D=1
M209 321 720 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=28380 $D=1
M210 318 314 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=23750 $D=1
M211 319 315 321 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=28380 $D=1
M212 320 43 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=23750 $D=1
M213 321 43 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=28380 $D=1
M214 242 44 320 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=23750 $D=1
M215 243 44 321 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=28380 $D=1
M216 322 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=23750 $D=1
M217 323 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=28380 $D=1
M218 6 45 324 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=23750 $D=1
M219 7 45 325 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=28380 $D=1
M220 326 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=23750 $D=1
M221 327 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=28380 $D=1
M222 328 45 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=23750 $D=1
M223 329 45 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=28380 $D=1
M224 6 328 721 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=23750 $D=1
M225 7 329 722 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=28380 $D=1
M226 330 721 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=23750 $D=1
M227 331 722 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=28380 $D=1
M228 328 324 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=23750 $D=1
M229 329 325 331 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=28380 $D=1
M230 330 46 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=23750 $D=1
M231 331 46 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=28380 $D=1
M232 242 47 330 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=23750 $D=1
M233 243 47 331 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=28380 $D=1
M234 332 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=23750 $D=1
M235 333 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=28380 $D=1
M236 6 48 334 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=23750 $D=1
M237 7 48 335 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=28380 $D=1
M238 336 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=23750 $D=1
M239 337 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=28380 $D=1
M240 338 48 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=23750 $D=1
M241 339 48 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=28380 $D=1
M242 6 338 723 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=23750 $D=1
M243 7 339 724 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=28380 $D=1
M244 340 723 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=23750 $D=1
M245 341 724 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=28380 $D=1
M246 338 334 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=23750 $D=1
M247 339 335 341 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=28380 $D=1
M248 340 49 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=23750 $D=1
M249 341 49 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=28380 $D=1
M250 242 50 340 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=23750 $D=1
M251 243 50 341 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=28380 $D=1
M252 342 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=23750 $D=1
M253 343 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=28380 $D=1
M254 6 51 344 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=23750 $D=1
M255 7 51 345 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=28380 $D=1
M256 346 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=23750 $D=1
M257 347 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=28380 $D=1
M258 348 51 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=23750 $D=1
M259 349 51 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=28380 $D=1
M260 6 348 725 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=23750 $D=1
M261 7 349 726 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=28380 $D=1
M262 350 725 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=23750 $D=1
M263 351 726 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=28380 $D=1
M264 348 344 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=23750 $D=1
M265 349 345 351 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=28380 $D=1
M266 350 52 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=23750 $D=1
M267 351 52 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=28380 $D=1
M268 242 53 350 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=23750 $D=1
M269 243 53 351 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=28380 $D=1
M270 352 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=23750 $D=1
M271 353 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=28380 $D=1
M272 6 54 354 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=23750 $D=1
M273 7 54 355 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=28380 $D=1
M274 356 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=23750 $D=1
M275 357 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=28380 $D=1
M276 358 54 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=23750 $D=1
M277 359 54 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=28380 $D=1
M278 6 358 727 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=23750 $D=1
M279 7 359 728 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=28380 $D=1
M280 360 727 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=23750 $D=1
M281 361 728 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=28380 $D=1
M282 358 354 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=23750 $D=1
M283 359 355 361 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=28380 $D=1
M284 360 55 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=23750 $D=1
M285 361 55 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=28380 $D=1
M286 242 56 360 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=23750 $D=1
M287 243 56 361 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=28380 $D=1
M288 362 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=23750 $D=1
M289 363 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=28380 $D=1
M290 6 57 364 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=23750 $D=1
M291 7 57 365 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=28380 $D=1
M292 366 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=23750 $D=1
M293 367 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=28380 $D=1
M294 368 57 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=23750 $D=1
M295 369 57 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=28380 $D=1
M296 6 368 729 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=23750 $D=1
M297 7 369 730 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=28380 $D=1
M298 370 729 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=23750 $D=1
M299 371 730 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=28380 $D=1
M300 368 364 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=23750 $D=1
M301 369 365 371 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=28380 $D=1
M302 370 58 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=23750 $D=1
M303 371 58 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=28380 $D=1
M304 242 59 370 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=23750 $D=1
M305 243 59 371 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=28380 $D=1
M306 372 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=23750 $D=1
M307 373 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=28380 $D=1
M308 6 60 374 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=23750 $D=1
M309 7 60 375 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=28380 $D=1
M310 376 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=23750 $D=1
M311 377 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=28380 $D=1
M312 378 60 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=23750 $D=1
M313 379 60 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=28380 $D=1
M314 6 378 731 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=23750 $D=1
M315 7 379 732 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=28380 $D=1
M316 380 731 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=23750 $D=1
M317 381 732 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=28380 $D=1
M318 378 374 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=23750 $D=1
M319 379 375 381 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=28380 $D=1
M320 380 61 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=23750 $D=1
M321 381 61 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=28380 $D=1
M322 242 62 380 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=23750 $D=1
M323 243 62 381 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=28380 $D=1
M324 382 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=23750 $D=1
M325 383 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=28380 $D=1
M326 6 63 384 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=23750 $D=1
M327 7 63 385 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=28380 $D=1
M328 386 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=23750 $D=1
M329 387 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=28380 $D=1
M330 388 63 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=23750 $D=1
M331 389 63 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=28380 $D=1
M332 6 388 733 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=23750 $D=1
M333 7 389 734 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=28380 $D=1
M334 390 733 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=23750 $D=1
M335 391 734 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=28380 $D=1
M336 388 384 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=23750 $D=1
M337 389 385 391 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=28380 $D=1
M338 390 64 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=23750 $D=1
M339 391 64 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=28380 $D=1
M340 242 65 390 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=23750 $D=1
M341 243 65 391 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=28380 $D=1
M342 392 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=23750 $D=1
M343 393 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=28380 $D=1
M344 6 66 394 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=23750 $D=1
M345 7 66 395 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=28380 $D=1
M346 396 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=23750 $D=1
M347 397 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=28380 $D=1
M348 398 66 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=23750 $D=1
M349 399 66 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=28380 $D=1
M350 6 398 735 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=23750 $D=1
M351 7 399 736 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=28380 $D=1
M352 400 735 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=23750 $D=1
M353 401 736 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=28380 $D=1
M354 398 394 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=23750 $D=1
M355 399 395 401 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=28380 $D=1
M356 400 67 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=23750 $D=1
M357 401 67 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=28380 $D=1
M358 242 68 400 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=23750 $D=1
M359 243 68 401 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=28380 $D=1
M360 402 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=23750 $D=1
M361 403 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=28380 $D=1
M362 6 69 404 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=23750 $D=1
M363 7 69 405 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=28380 $D=1
M364 406 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=23750 $D=1
M365 407 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=28380 $D=1
M366 408 69 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=23750 $D=1
M367 409 69 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=28380 $D=1
M368 6 408 737 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=23750 $D=1
M369 7 409 738 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=28380 $D=1
M370 410 737 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=23750 $D=1
M371 411 738 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=28380 $D=1
M372 408 404 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=23750 $D=1
M373 409 405 411 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=28380 $D=1
M374 410 70 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=23750 $D=1
M375 411 70 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=28380 $D=1
M376 242 71 410 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=23750 $D=1
M377 243 71 411 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=28380 $D=1
M378 412 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=23750 $D=1
M379 413 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=28380 $D=1
M380 6 72 414 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=23750 $D=1
M381 7 72 415 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=28380 $D=1
M382 416 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=23750 $D=1
M383 417 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=28380 $D=1
M384 418 72 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=23750 $D=1
M385 419 72 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=28380 $D=1
M386 6 418 739 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=23750 $D=1
M387 7 419 740 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=28380 $D=1
M388 420 739 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=23750 $D=1
M389 421 740 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=28380 $D=1
M390 418 414 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=23750 $D=1
M391 419 415 421 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=28380 $D=1
M392 420 73 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=23750 $D=1
M393 421 73 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=28380 $D=1
M394 242 74 420 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=23750 $D=1
M395 243 74 421 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=28380 $D=1
M396 422 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=23750 $D=1
M397 423 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=28380 $D=1
M398 6 75 424 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=23750 $D=1
M399 7 75 425 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=28380 $D=1
M400 426 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=23750 $D=1
M401 427 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=28380 $D=1
M402 428 75 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=23750 $D=1
M403 429 75 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=28380 $D=1
M404 6 428 741 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=23750 $D=1
M405 7 429 742 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=28380 $D=1
M406 430 741 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=23750 $D=1
M407 431 742 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=28380 $D=1
M408 428 424 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=23750 $D=1
M409 429 425 431 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=28380 $D=1
M410 430 76 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=23750 $D=1
M411 431 76 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=28380 $D=1
M412 242 77 430 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=23750 $D=1
M413 243 77 431 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=28380 $D=1
M414 432 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=23750 $D=1
M415 433 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=28380 $D=1
M416 6 78 434 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=23750 $D=1
M417 7 78 435 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=28380 $D=1
M418 436 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=23750 $D=1
M419 437 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=28380 $D=1
M420 438 78 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=23750 $D=1
M421 439 78 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=28380 $D=1
M422 6 438 743 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=23750 $D=1
M423 7 439 744 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=28380 $D=1
M424 440 743 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=23750 $D=1
M425 441 744 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=28380 $D=1
M426 438 434 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=23750 $D=1
M427 439 435 441 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=28380 $D=1
M428 440 79 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=23750 $D=1
M429 441 79 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=28380 $D=1
M430 242 80 440 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=23750 $D=1
M431 243 80 441 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=28380 $D=1
M432 442 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=23750 $D=1
M433 443 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=28380 $D=1
M434 6 81 444 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=23750 $D=1
M435 7 81 445 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=28380 $D=1
M436 446 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=23750 $D=1
M437 447 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=28380 $D=1
M438 448 81 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=23750 $D=1
M439 449 81 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=28380 $D=1
M440 6 448 745 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=23750 $D=1
M441 7 449 746 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=28380 $D=1
M442 450 745 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=23750 $D=1
M443 451 746 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=28380 $D=1
M444 448 444 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=23750 $D=1
M445 449 445 451 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=28380 $D=1
M446 450 82 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=23750 $D=1
M447 451 82 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=28380 $D=1
M448 242 83 450 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=23750 $D=1
M449 243 83 451 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=28380 $D=1
M450 452 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=23750 $D=1
M451 453 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=28380 $D=1
M452 6 84 454 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=23750 $D=1
M453 7 84 455 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=28380 $D=1
M454 456 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=23750 $D=1
M455 457 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=28380 $D=1
M456 458 84 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=23750 $D=1
M457 459 84 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=28380 $D=1
M458 6 458 747 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=23750 $D=1
M459 7 459 748 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=28380 $D=1
M460 460 747 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=23750 $D=1
M461 461 748 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=28380 $D=1
M462 458 454 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=23750 $D=1
M463 459 455 461 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=28380 $D=1
M464 460 85 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=23750 $D=1
M465 461 85 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=28380 $D=1
M466 242 86 460 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=23750 $D=1
M467 243 86 461 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=28380 $D=1
M468 462 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=23750 $D=1
M469 463 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=28380 $D=1
M470 6 87 464 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=23750 $D=1
M471 7 87 465 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=28380 $D=1
M472 466 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=23750 $D=1
M473 467 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=28380 $D=1
M474 468 87 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=23750 $D=1
M475 469 87 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=28380 $D=1
M476 6 468 749 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=23750 $D=1
M477 7 469 750 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=28380 $D=1
M478 470 749 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=23750 $D=1
M479 471 750 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=28380 $D=1
M480 468 464 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=23750 $D=1
M481 469 465 471 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=28380 $D=1
M482 470 88 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=23750 $D=1
M483 471 88 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=28380 $D=1
M484 242 89 470 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=23750 $D=1
M485 243 89 471 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=28380 $D=1
M486 472 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=23750 $D=1
M487 473 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=28380 $D=1
M488 6 90 474 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=23750 $D=1
M489 7 90 475 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=28380 $D=1
M490 476 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=23750 $D=1
M491 477 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=28380 $D=1
M492 478 90 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=23750 $D=1
M493 479 90 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=28380 $D=1
M494 6 478 751 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=23750 $D=1
M495 7 479 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=28380 $D=1
M496 480 751 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=23750 $D=1
M497 481 752 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=28380 $D=1
M498 478 474 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=23750 $D=1
M499 479 475 481 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=28380 $D=1
M500 480 91 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=23750 $D=1
M501 481 91 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=28380 $D=1
M502 242 92 480 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=23750 $D=1
M503 243 92 481 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=28380 $D=1
M504 482 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=23750 $D=1
M505 483 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=28380 $D=1
M506 6 93 484 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=23750 $D=1
M507 7 93 485 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=28380 $D=1
M508 486 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=23750 $D=1
M509 487 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=28380 $D=1
M510 488 93 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=23750 $D=1
M511 489 93 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=28380 $D=1
M512 6 488 753 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=23750 $D=1
M513 7 489 754 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=28380 $D=1
M514 490 753 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=23750 $D=1
M515 491 754 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=28380 $D=1
M516 488 484 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=23750 $D=1
M517 489 485 491 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=28380 $D=1
M518 490 94 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=23750 $D=1
M519 491 94 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=28380 $D=1
M520 242 95 490 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=23750 $D=1
M521 243 95 491 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=28380 $D=1
M522 492 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=23750 $D=1
M523 493 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=28380 $D=1
M524 6 96 494 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=23750 $D=1
M525 7 96 495 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=28380 $D=1
M526 496 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=23750 $D=1
M527 497 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=28380 $D=1
M528 498 96 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=23750 $D=1
M529 499 96 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=28380 $D=1
M530 6 498 755 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=23750 $D=1
M531 7 499 756 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=28380 $D=1
M532 500 755 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=23750 $D=1
M533 501 756 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=28380 $D=1
M534 498 494 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=23750 $D=1
M535 499 495 501 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=28380 $D=1
M536 500 97 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=23750 $D=1
M537 501 97 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=28380 $D=1
M538 242 98 500 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=23750 $D=1
M539 243 98 501 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=28380 $D=1
M540 502 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=23750 $D=1
M541 503 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=28380 $D=1
M542 6 99 504 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=23750 $D=1
M543 7 99 505 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=28380 $D=1
M544 506 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=23750 $D=1
M545 507 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=28380 $D=1
M546 508 99 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=23750 $D=1
M547 509 99 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=28380 $D=1
M548 6 508 757 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=23750 $D=1
M549 7 509 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=28380 $D=1
M550 510 757 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=23750 $D=1
M551 511 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=28380 $D=1
M552 508 504 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=23750 $D=1
M553 509 505 511 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=28380 $D=1
M554 510 100 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=23750 $D=1
M555 511 100 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=28380 $D=1
M556 242 101 510 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=23750 $D=1
M557 243 101 511 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=28380 $D=1
M558 512 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=23750 $D=1
M559 513 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=28380 $D=1
M560 6 102 514 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=23750 $D=1
M561 7 102 515 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=28380 $D=1
M562 516 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=23750 $D=1
M563 517 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=28380 $D=1
M564 518 102 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=23750 $D=1
M565 519 102 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=28380 $D=1
M566 6 518 759 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=23750 $D=1
M567 7 519 760 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=28380 $D=1
M568 520 759 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=23750 $D=1
M569 521 760 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=28380 $D=1
M570 518 514 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=23750 $D=1
M571 519 515 521 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=28380 $D=1
M572 520 103 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=23750 $D=1
M573 521 103 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=28380 $D=1
M574 242 104 520 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=23750 $D=1
M575 243 104 521 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=28380 $D=1
M576 522 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=23750 $D=1
M577 523 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=28380 $D=1
M578 6 105 524 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=23750 $D=1
M579 7 105 525 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=28380 $D=1
M580 526 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=23750 $D=1
M581 527 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=28380 $D=1
M582 528 105 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=23750 $D=1
M583 529 105 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=28380 $D=1
M584 6 528 761 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=23750 $D=1
M585 7 529 762 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=28380 $D=1
M586 530 761 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=23750 $D=1
M587 531 762 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=28380 $D=1
M588 528 524 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=23750 $D=1
M589 529 525 531 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=28380 $D=1
M590 530 106 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=23750 $D=1
M591 531 106 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=28380 $D=1
M592 242 108 530 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=23750 $D=1
M593 243 108 531 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=28380 $D=1
M594 532 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=23750 $D=1
M595 533 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=28380 $D=1
M596 6 109 534 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=23750 $D=1
M597 7 109 535 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=28380 $D=1
M598 536 110 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=23750 $D=1
M599 537 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=28380 $D=1
M600 538 109 228 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=23750 $D=1
M601 539 109 229 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=28380 $D=1
M602 6 538 763 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=23750 $D=1
M603 7 539 764 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=28380 $D=1
M604 540 763 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=23750 $D=1
M605 541 764 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=28380 $D=1
M606 538 534 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=23750 $D=1
M607 539 535 541 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=28380 $D=1
M608 540 110 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=23750 $D=1
M609 541 110 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=28380 $D=1
M610 242 112 540 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=23750 $D=1
M611 243 112 541 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=28380 $D=1
M612 542 112 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=23750 $D=1
M613 543 112 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=28380 $D=1
M614 6 113 544 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=23750 $D=1
M615 7 113 545 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=28380 $D=1
M616 546 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=23750 $D=1
M617 547 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=28380 $D=1
M618 6 114 238 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=23750 $D=1
M619 7 114 239 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=28380 $D=1
M620 242 113 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=23750 $D=1
M621 243 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=28380 $D=1
M622 6 550 548 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=23750 $D=1
M623 7 551 549 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=28380 $D=1
M624 550 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=23750 $D=1
M625 551 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=28380 $D=1
M626 765 238 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=23750 $D=1
M627 766 239 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=28380 $D=1
M628 552 548 765 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=23750 $D=1
M629 553 549 766 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=28380 $D=1
M630 6 552 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=23750 $D=1
M631 7 553 555 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=28380 $D=1
M632 767 554 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=23750 $D=1
M633 768 555 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=28380 $D=1
M634 552 550 767 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=23750 $D=1
M635 553 551 768 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=28380 $D=1
M636 6 558 556 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=23750 $D=1
M637 7 559 557 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=28380 $D=1
M638 558 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=23750 $D=1
M639 559 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=28380 $D=1
M640 769 242 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=23750 $D=1
M641 770 243 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=28380 $D=1
M642 560 556 769 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=23750 $D=1
M643 561 557 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=28380 $D=1
M644 6 560 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=23750 $D=1
M645 7 561 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=28380 $D=1
M646 771 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=23750 $D=1
M647 772 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=28380 $D=1
M648 560 558 771 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=23750 $D=1
M649 561 559 772 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=28380 $D=1
M650 562 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=23750 $D=1
M651 563 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=28380 $D=1
M652 564 562 554 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=23750 $D=1
M653 565 563 555 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=28380 $D=1
M654 121 120 564 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=23750 $D=1
M655 122 120 565 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=28380 $D=1
M656 566 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=23750 $D=1
M657 567 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=28380 $D=1
M658 568 566 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=23750 $D=1
M659 569 567 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=28380 $D=1
M660 773 123 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=23750 $D=1
M661 774 123 569 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=28380 $D=1
M662 6 118 773 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=23750 $D=1
M663 7 119 774 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=28380 $D=1
M664 570 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=23750 $D=1
M665 571 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=28380 $D=1
M666 572 570 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=23750 $D=1
M667 573 571 569 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=28380 $D=1
M668 12 124 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=23750 $D=1
M669 13 124 573 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=28380 $D=1
M670 576 574 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=23750 $D=1
M671 577 575 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=28380 $D=1
M672 6 580 578 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=23750 $D=1
M673 7 581 579 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=28380 $D=1
M674 582 564 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=23750 $D=1
M675 583 565 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=28380 $D=1
M676 580 582 574 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=23750 $D=1
M677 581 583 575 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=28380 $D=1
M678 576 564 580 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=23750 $D=1
M679 577 565 581 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=28380 $D=1
M680 584 578 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=23750 $D=1
M681 585 579 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=28380 $D=1
M682 125 584 572 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=23750 $D=1
M683 574 585 573 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=28380 $D=1
M684 564 578 125 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=23750 $D=1
M685 565 579 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=28380 $D=1
M686 586 125 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=23750 $D=1
M687 587 574 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=28380 $D=1
M688 588 578 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=23750 $D=1
M689 589 579 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=28380 $D=1
M690 590 588 586 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=23750 $D=1
M691 591 589 587 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=28380 $D=1
M692 572 578 590 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=23750 $D=1
M693 573 579 591 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=28380 $D=1
M694 592 564 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=23750 $D=1
M695 593 565 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=28380 $D=1
M696 6 572 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=23750 $D=1
M697 7 573 593 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=28380 $D=1
M698 594 590 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=23750 $D=1
M699 595 591 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=28380 $D=1
M700 793 564 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=23750 $D=1
M701 794 565 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=28380 $D=1
M702 596 572 793 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=23750 $D=1
M703 597 573 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=28380 $D=1
M704 795 564 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=23750 $D=1
M705 796 565 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=28380 $D=1
M706 598 572 795 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=23750 $D=1
M707 599 573 796 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=28380 $D=1
M708 602 564 600 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=23750 $D=1
M709 603 565 601 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=28380 $D=1
M710 600 572 602 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=23750 $D=1
M711 601 573 603 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=28380 $D=1
M712 6 598 600 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=23750 $D=1
M713 7 599 601 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=28380 $D=1
M714 604 128 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=23750 $D=1
M715 605 128 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=28380 $D=1
M716 606 604 592 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=23750 $D=1
M717 607 605 593 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=28380 $D=1
M718 596 128 606 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=23750 $D=1
M719 597 128 607 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=28380 $D=1
M720 608 604 594 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=23750 $D=1
M721 609 605 595 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=28380 $D=1
M722 602 128 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=23750 $D=1
M723 603 128 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=28380 $D=1
M724 610 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=23750 $D=1
M725 611 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=28380 $D=1
M726 612 610 608 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=23750 $D=1
M727 613 611 609 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=28380 $D=1
M728 606 129 612 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=23750 $D=1
M729 607 129 613 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=28380 $D=1
M730 14 612 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=23750 $D=1
M731 15 613 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=28380 $D=1
M732 614 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=23750 $D=1
M733 615 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=28380 $D=1
M734 616 614 131 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=23750 $D=1
M735 617 615 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=28380 $D=1
M736 133 130 616 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=23750 $D=1
M737 134 130 617 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=28380 $D=1
M738 618 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=23750 $D=1
M739 619 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=28380 $D=1
M740 620 618 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=23750 $D=1
M741 621 619 136 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=28380 $D=1
M742 137 130 620 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=23750 $D=1
M743 138 130 621 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=28380 $D=1
M744 622 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=23750 $D=1
M745 623 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=28380 $D=1
M746 624 622 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=23750 $D=1
M747 625 623 126 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=28380 $D=1
M748 139 130 624 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=23750 $D=1
M749 140 130 625 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=28380 $D=1
M750 626 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=23750 $D=1
M751 627 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=28380 $D=1
M752 628 626 142 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=23750 $D=1
M753 629 627 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=28380 $D=1
M754 144 130 628 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=23750 $D=1
M755 144 130 629 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=28380 $D=1
M756 630 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=23750 $D=1
M757 631 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=28380 $D=1
M758 632 630 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=23750 $D=1
M759 633 631 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=28380 $D=1
M760 144 130 632 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=23750 $D=1
M761 144 130 633 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=28380 $D=1
M762 6 564 775 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=23750 $D=1
M763 7 565 776 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=28380 $D=1
M764 134 775 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=23750 $D=1
M765 131 776 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=28380 $D=1
M766 634 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=23750 $D=1
M767 635 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=28380 $D=1
M768 148 634 134 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=23750 $D=1
M769 149 635 131 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=28380 $D=1
M770 616 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=23750 $D=1
M771 617 147 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=28380 $D=1
M772 636 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=23750 $D=1
M773 637 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=28380 $D=1
M774 151 636 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=23750 $D=1
M775 107 637 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=28380 $D=1
M776 620 150 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=23750 $D=1
M777 621 150 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=28380 $D=1
M778 638 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=23750 $D=1
M779 639 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=28380 $D=1
M780 153 638 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=23750 $D=1
M781 115 639 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=28380 $D=1
M782 624 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=23750 $D=1
M783 625 152 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=28380 $D=1
M784 640 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=23750 $D=1
M785 641 154 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=28380 $D=1
M786 155 640 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=23750 $D=1
M787 156 641 115 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=28380 $D=1
M788 628 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=23750 $D=1
M789 629 154 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=28380 $D=1
M790 642 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=23750 $D=1
M791 643 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=28380 $D=1
M792 214 642 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=23750 $D=1
M793 215 643 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=28380 $D=1
M794 632 157 214 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=23750 $D=1
M795 633 157 215 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=28380 $D=1
M796 644 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=23750 $D=1
M797 645 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=28380 $D=1
M798 646 644 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=23750 $D=1
M799 647 645 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=28380 $D=1
M800 12 158 646 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=23750 $D=1
M801 13 158 647 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=28380 $D=1
M802 797 554 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=23750 $D=1
M803 798 555 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=28380 $D=1
M804 648 646 797 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=23750 $D=1
M805 649 647 798 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=28380 $D=1
M806 652 554 650 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=23750 $D=1
M807 653 555 651 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=28380 $D=1
M808 650 646 652 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=23750 $D=1
M809 651 647 653 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=28380 $D=1
M810 6 648 650 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=23750 $D=1
M811 7 649 651 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=28380 $D=1
M812 799 159 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=23750 $D=1
M813 800 654 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=28380 $D=1
M814 777 652 799 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=23750 $D=1
M815 778 653 800 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=28380 $D=1
M816 654 777 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=23750 $D=1
M817 160 778 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=28380 $D=1
M818 655 554 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=23750 $D=1
M819 656 555 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=28380 $D=1
M820 6 657 655 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=23750 $D=1
M821 7 658 656 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=28380 $D=1
M822 657 646 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=23750 $D=1
M823 658 647 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=28380 $D=1
M824 801 655 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=23750 $D=1
M825 802 656 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=28380 $D=1
M826 659 159 801 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=23750 $D=1
M827 660 654 802 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=28380 $D=1
M828 662 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=23750 $D=1
M829 663 661 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=28380 $D=1
M830 803 659 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=23750 $D=1
M831 804 660 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=28380 $D=1
M832 661 662 803 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=23750 $D=1
M833 162 663 804 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=28380 $D=1
M834 665 664 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=23750 $D=1
M835 666 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=28380 $D=1
M836 6 669 667 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=23750 $D=1
M837 7 670 668 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=28380 $D=1
M838 671 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=23750 $D=1
M839 672 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=28380 $D=1
M840 669 671 664 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=23750 $D=1
M841 670 672 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=28380 $D=1
M842 665 121 669 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=23750 $D=1
M843 666 122 670 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=28380 $D=1
M844 673 667 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=23750 $D=1
M845 674 668 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=28380 $D=1
M846 164 673 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=23750 $D=1
M847 664 674 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=28380 $D=1
M848 121 667 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=23750 $D=1
M849 122 668 664 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=28380 $D=1
M850 675 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=23750 $D=1
M851 676 664 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=28380 $D=1
M852 677 667 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=23750 $D=1
M853 678 668 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=28380 $D=1
M854 216 677 675 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=23750 $D=1
M855 217 678 676 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=28380 $D=1
M856 6 667 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=23750 $D=1
M857 7 668 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=28380 $D=1
M858 679 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=23750 $D=1
M859 680 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=28380 $D=1
M860 681 679 216 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=23750 $D=1
M861 682 680 217 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=28380 $D=1
M862 14 165 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=23750 $D=1
M863 15 165 682 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=28380 $D=1
M864 683 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=23750 $D=1
M865 684 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=28380 $D=1
M866 166 683 681 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=23750 $D=1
M867 166 684 682 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=28380 $D=1
M868 6 166 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=23750 $D=1
M869 7 166 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=28380 $D=1
M870 685 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=23750 $D=1
M871 686 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=28380 $D=1
M872 6 685 687 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=23750 $D=1
M873 7 686 688 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=28380 $D=1
M874 689 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=23750 $D=1
M875 690 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=28380 $D=1
M876 691 685 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=23750 $D=1
M877 692 686 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=28380 $D=1
M878 6 691 779 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=23750 $D=1
M879 7 692 780 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=28380 $D=1
M880 693 779 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=23750 $D=1
M881 694 780 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=28380 $D=1
M882 691 687 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=23750 $D=1
M883 692 688 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=28380 $D=1
M884 695 116 693 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=23750 $D=1
M885 696 116 694 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=28380 $D=1
M886 6 699 697 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=23750 $D=1
M887 7 700 698 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=28380 $D=1
M888 699 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=23750 $D=1
M889 700 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=28380 $D=1
M890 781 695 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=23750 $D=1
M891 782 696 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=28380 $D=1
M892 701 697 781 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=23750 $D=1
M893 702 698 782 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=28380 $D=1
M894 6 701 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=23750 $D=1
M895 7 702 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=28380 $D=1
M896 783 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=23750 $D=1
M897 784 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=28380 $D=1
M898 701 699 783 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=23750 $D=1
M899 702 700 784 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=28380 $D=1
M900 190 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=25000 $D=0
M901 191 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=29630 $D=0
M902 192 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=25000 $D=0
M903 193 1 3 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=29630 $D=0
M904 6 190 192 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=25000 $D=0
M905 7 191 193 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=29630 $D=0
M906 194 1 4 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=25000 $D=0
M907 195 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=29630 $D=0
M908 5 190 194 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=25000 $D=0
M909 5 191 195 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=29630 $D=0
M910 196 1 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=25000 $D=0
M911 197 1 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=29630 $D=0
M912 6 190 196 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=25000 $D=0
M913 7 191 197 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=29630 $D=0
M914 200 9 196 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=25000 $D=0
M915 201 9 197 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=29630 $D=0
M916 198 9 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=25000 $D=0
M917 199 9 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=29630 $D=0
M918 202 9 194 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=25000 $D=0
M919 203 9 195 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=29630 $D=0
M920 192 198 202 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=25000 $D=0
M921 193 199 203 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=29630 $D=0
M922 204 10 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=25000 $D=0
M923 205 10 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=29630 $D=0
M924 206 10 202 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=25000 $D=0
M925 207 10 203 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=29630 $D=0
M926 200 204 206 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=25000 $D=0
M927 201 205 207 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=29630 $D=0
M928 208 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=25000 $D=0
M929 209 11 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=29630 $D=0
M930 210 11 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=25000 $D=0
M931 211 11 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=29630 $D=0
M932 12 208 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=25000 $D=0
M933 13 209 211 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=29630 $D=0
M934 212 11 14 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=25000 $D=0
M935 213 11 15 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=29630 $D=0
M936 214 208 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=25000 $D=0
M937 215 209 213 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=29630 $D=0
M938 218 11 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=25000 $D=0
M939 219 11 217 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=29630 $D=0
M940 206 208 218 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=25000 $D=0
M941 207 209 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=29630 $D=0
M942 222 16 218 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=25000 $D=0
M943 223 16 219 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=29630 $D=0
M944 220 16 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=25000 $D=0
M945 221 16 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=29630 $D=0
M946 224 16 212 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=25000 $D=0
M947 225 16 213 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=29630 $D=0
M948 210 220 224 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=25000 $D=0
M949 211 221 225 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=29630 $D=0
M950 226 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=25000 $D=0
M951 227 17 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=29630 $D=0
M952 228 17 224 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=25000 $D=0
M953 229 17 225 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=29630 $D=0
M954 222 226 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=25000 $D=0
M955 223 227 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=29630 $D=0
M956 167 18 230 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=25000 $D=0
M957 168 18 231 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=29630 $D=0
M958 232 19 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=25000 $D=0
M959 233 19 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=29630 $D=0
M960 234 230 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=25000 $D=0
M961 235 231 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=29630 $D=0
M962 167 234 703 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=25000 $D=0
M963 168 235 704 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=29630 $D=0
M964 236 703 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=25000 $D=0
M965 237 704 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=29630 $D=0
M966 234 18 236 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=25000 $D=0
M967 235 18 237 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=29630 $D=0
M968 236 232 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=25000 $D=0
M969 237 233 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=29630 $D=0
M970 242 240 236 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=25000 $D=0
M971 243 241 237 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=29630 $D=0
M972 240 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=25000 $D=0
M973 241 20 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=29630 $D=0
M974 167 21 244 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=25000 $D=0
M975 168 21 245 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=29630 $D=0
M976 246 22 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=25000 $D=0
M977 247 22 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=29630 $D=0
M978 248 244 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=25000 $D=0
M979 249 245 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=29630 $D=0
M980 167 248 705 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=25000 $D=0
M981 168 249 706 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=29630 $D=0
M982 250 705 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=25000 $D=0
M983 251 706 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=29630 $D=0
M984 248 21 250 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=25000 $D=0
M985 249 21 251 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=29630 $D=0
M986 250 246 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=25000 $D=0
M987 251 247 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=29630 $D=0
M988 242 252 250 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=25000 $D=0
M989 243 253 251 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=29630 $D=0
M990 252 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=25000 $D=0
M991 253 23 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=29630 $D=0
M992 167 24 254 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=25000 $D=0
M993 168 24 255 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=29630 $D=0
M994 256 25 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=25000 $D=0
M995 257 25 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=29630 $D=0
M996 258 254 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=25000 $D=0
M997 259 255 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=29630 $D=0
M998 167 258 707 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=25000 $D=0
M999 168 259 708 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=29630 $D=0
M1000 260 707 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=25000 $D=0
M1001 261 708 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=29630 $D=0
M1002 258 24 260 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=25000 $D=0
M1003 259 24 261 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=29630 $D=0
M1004 260 256 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=25000 $D=0
M1005 261 257 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=29630 $D=0
M1006 242 262 260 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=25000 $D=0
M1007 243 263 261 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=29630 $D=0
M1008 262 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=25000 $D=0
M1009 263 26 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=29630 $D=0
M1010 167 27 264 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=25000 $D=0
M1011 168 27 265 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=29630 $D=0
M1012 266 28 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=25000 $D=0
M1013 267 28 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=29630 $D=0
M1014 268 264 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=25000 $D=0
M1015 269 265 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=29630 $D=0
M1016 167 268 709 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=25000 $D=0
M1017 168 269 710 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=29630 $D=0
M1018 270 709 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=25000 $D=0
M1019 271 710 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=29630 $D=0
M1020 268 27 270 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=25000 $D=0
M1021 269 27 271 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=29630 $D=0
M1022 270 266 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=25000 $D=0
M1023 271 267 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=29630 $D=0
M1024 242 272 270 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=25000 $D=0
M1025 243 273 271 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=29630 $D=0
M1026 272 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=25000 $D=0
M1027 273 29 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=29630 $D=0
M1028 167 30 274 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=25000 $D=0
M1029 168 30 275 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=29630 $D=0
M1030 276 31 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=25000 $D=0
M1031 277 31 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=29630 $D=0
M1032 278 274 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=25000 $D=0
M1033 279 275 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=29630 $D=0
M1034 167 278 711 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=25000 $D=0
M1035 168 279 712 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=29630 $D=0
M1036 280 711 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=25000 $D=0
M1037 281 712 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=29630 $D=0
M1038 278 30 280 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=25000 $D=0
M1039 279 30 281 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=29630 $D=0
M1040 280 276 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=25000 $D=0
M1041 281 277 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=29630 $D=0
M1042 242 282 280 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=25000 $D=0
M1043 243 283 281 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=29630 $D=0
M1044 282 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=25000 $D=0
M1045 283 32 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=29630 $D=0
M1046 167 33 284 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=25000 $D=0
M1047 168 33 285 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=29630 $D=0
M1048 286 34 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=25000 $D=0
M1049 287 34 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=29630 $D=0
M1050 288 284 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=25000 $D=0
M1051 289 285 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=29630 $D=0
M1052 167 288 713 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=25000 $D=0
M1053 168 289 714 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=29630 $D=0
M1054 290 713 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=25000 $D=0
M1055 291 714 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=29630 $D=0
M1056 288 33 290 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=25000 $D=0
M1057 289 33 291 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=29630 $D=0
M1058 290 286 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=25000 $D=0
M1059 291 287 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=29630 $D=0
M1060 242 292 290 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=25000 $D=0
M1061 243 293 291 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=29630 $D=0
M1062 292 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=25000 $D=0
M1063 293 35 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=29630 $D=0
M1064 167 36 294 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=25000 $D=0
M1065 168 36 295 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=29630 $D=0
M1066 296 37 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=25000 $D=0
M1067 297 37 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=29630 $D=0
M1068 298 294 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=25000 $D=0
M1069 299 295 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=29630 $D=0
M1070 167 298 715 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=25000 $D=0
M1071 168 299 716 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=29630 $D=0
M1072 300 715 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=25000 $D=0
M1073 301 716 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=29630 $D=0
M1074 298 36 300 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=25000 $D=0
M1075 299 36 301 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=29630 $D=0
M1076 300 296 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=25000 $D=0
M1077 301 297 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=29630 $D=0
M1078 242 302 300 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=25000 $D=0
M1079 243 303 301 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=29630 $D=0
M1080 302 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=25000 $D=0
M1081 303 38 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=29630 $D=0
M1082 167 39 304 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=25000 $D=0
M1083 168 39 305 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=29630 $D=0
M1084 306 40 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=25000 $D=0
M1085 307 40 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=29630 $D=0
M1086 308 304 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=25000 $D=0
M1087 309 305 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=29630 $D=0
M1088 167 308 717 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=25000 $D=0
M1089 168 309 718 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=29630 $D=0
M1090 310 717 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=25000 $D=0
M1091 311 718 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=29630 $D=0
M1092 308 39 310 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=25000 $D=0
M1093 309 39 311 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=29630 $D=0
M1094 310 306 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=25000 $D=0
M1095 311 307 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=29630 $D=0
M1096 242 312 310 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=25000 $D=0
M1097 243 313 311 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=29630 $D=0
M1098 312 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=25000 $D=0
M1099 313 41 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=29630 $D=0
M1100 167 42 314 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=25000 $D=0
M1101 168 42 315 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=29630 $D=0
M1102 316 43 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=25000 $D=0
M1103 317 43 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=29630 $D=0
M1104 318 314 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=25000 $D=0
M1105 319 315 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=29630 $D=0
M1106 167 318 719 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=25000 $D=0
M1107 168 319 720 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=29630 $D=0
M1108 320 719 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=25000 $D=0
M1109 321 720 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=29630 $D=0
M1110 318 42 320 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=25000 $D=0
M1111 319 42 321 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=29630 $D=0
M1112 320 316 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=25000 $D=0
M1113 321 317 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=29630 $D=0
M1114 242 322 320 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=25000 $D=0
M1115 243 323 321 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=29630 $D=0
M1116 322 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=25000 $D=0
M1117 323 44 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=29630 $D=0
M1118 167 45 324 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=25000 $D=0
M1119 168 45 325 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=29630 $D=0
M1120 326 46 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=25000 $D=0
M1121 327 46 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=29630 $D=0
M1122 328 324 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=25000 $D=0
M1123 329 325 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=29630 $D=0
M1124 167 328 721 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=25000 $D=0
M1125 168 329 722 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=29630 $D=0
M1126 330 721 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=25000 $D=0
M1127 331 722 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=29630 $D=0
M1128 328 45 330 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=25000 $D=0
M1129 329 45 331 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=29630 $D=0
M1130 330 326 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=25000 $D=0
M1131 331 327 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=29630 $D=0
M1132 242 332 330 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=25000 $D=0
M1133 243 333 331 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=29630 $D=0
M1134 332 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=25000 $D=0
M1135 333 47 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=29630 $D=0
M1136 167 48 334 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=25000 $D=0
M1137 168 48 335 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=29630 $D=0
M1138 336 49 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=25000 $D=0
M1139 337 49 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=29630 $D=0
M1140 338 334 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=25000 $D=0
M1141 339 335 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=29630 $D=0
M1142 167 338 723 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=25000 $D=0
M1143 168 339 724 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=29630 $D=0
M1144 340 723 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=25000 $D=0
M1145 341 724 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=29630 $D=0
M1146 338 48 340 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=25000 $D=0
M1147 339 48 341 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=29630 $D=0
M1148 340 336 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=25000 $D=0
M1149 341 337 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=29630 $D=0
M1150 242 342 340 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=25000 $D=0
M1151 243 343 341 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=29630 $D=0
M1152 342 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=25000 $D=0
M1153 343 50 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=29630 $D=0
M1154 167 51 344 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=25000 $D=0
M1155 168 51 345 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=29630 $D=0
M1156 346 52 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=25000 $D=0
M1157 347 52 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=29630 $D=0
M1158 348 344 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=25000 $D=0
M1159 349 345 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=29630 $D=0
M1160 167 348 725 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=25000 $D=0
M1161 168 349 726 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=29630 $D=0
M1162 350 725 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=25000 $D=0
M1163 351 726 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=29630 $D=0
M1164 348 51 350 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=25000 $D=0
M1165 349 51 351 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=29630 $D=0
M1166 350 346 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=25000 $D=0
M1167 351 347 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=29630 $D=0
M1168 242 352 350 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=25000 $D=0
M1169 243 353 351 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=29630 $D=0
M1170 352 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=25000 $D=0
M1171 353 53 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=29630 $D=0
M1172 167 54 354 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=25000 $D=0
M1173 168 54 355 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=29630 $D=0
M1174 356 55 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=25000 $D=0
M1175 357 55 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=29630 $D=0
M1176 358 354 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=25000 $D=0
M1177 359 355 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=29630 $D=0
M1178 167 358 727 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=25000 $D=0
M1179 168 359 728 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=29630 $D=0
M1180 360 727 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=25000 $D=0
M1181 361 728 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=29630 $D=0
M1182 358 54 360 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=25000 $D=0
M1183 359 54 361 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=29630 $D=0
M1184 360 356 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=25000 $D=0
M1185 361 357 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=29630 $D=0
M1186 242 362 360 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=25000 $D=0
M1187 243 363 361 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=29630 $D=0
M1188 362 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=25000 $D=0
M1189 363 56 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=29630 $D=0
M1190 167 57 364 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=25000 $D=0
M1191 168 57 365 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=29630 $D=0
M1192 366 58 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=25000 $D=0
M1193 367 58 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=29630 $D=0
M1194 368 364 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=25000 $D=0
M1195 369 365 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=29630 $D=0
M1196 167 368 729 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=25000 $D=0
M1197 168 369 730 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=29630 $D=0
M1198 370 729 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=25000 $D=0
M1199 371 730 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=29630 $D=0
M1200 368 57 370 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=25000 $D=0
M1201 369 57 371 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=29630 $D=0
M1202 370 366 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=25000 $D=0
M1203 371 367 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=29630 $D=0
M1204 242 372 370 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=25000 $D=0
M1205 243 373 371 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=29630 $D=0
M1206 372 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=25000 $D=0
M1207 373 59 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=29630 $D=0
M1208 167 60 374 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=25000 $D=0
M1209 168 60 375 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=29630 $D=0
M1210 376 61 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=25000 $D=0
M1211 377 61 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=29630 $D=0
M1212 378 374 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=25000 $D=0
M1213 379 375 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=29630 $D=0
M1214 167 378 731 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=25000 $D=0
M1215 168 379 732 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=29630 $D=0
M1216 380 731 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=25000 $D=0
M1217 381 732 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=29630 $D=0
M1218 378 60 380 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=25000 $D=0
M1219 379 60 381 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=29630 $D=0
M1220 380 376 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=25000 $D=0
M1221 381 377 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=29630 $D=0
M1222 242 382 380 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=25000 $D=0
M1223 243 383 381 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=29630 $D=0
M1224 382 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=25000 $D=0
M1225 383 62 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=29630 $D=0
M1226 167 63 384 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=25000 $D=0
M1227 168 63 385 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=29630 $D=0
M1228 386 64 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=25000 $D=0
M1229 387 64 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=29630 $D=0
M1230 388 384 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=25000 $D=0
M1231 389 385 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=29630 $D=0
M1232 167 388 733 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=25000 $D=0
M1233 168 389 734 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=29630 $D=0
M1234 390 733 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=25000 $D=0
M1235 391 734 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=29630 $D=0
M1236 388 63 390 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=25000 $D=0
M1237 389 63 391 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=29630 $D=0
M1238 390 386 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=25000 $D=0
M1239 391 387 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=29630 $D=0
M1240 242 392 390 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=25000 $D=0
M1241 243 393 391 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=29630 $D=0
M1242 392 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=25000 $D=0
M1243 393 65 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=29630 $D=0
M1244 167 66 394 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=25000 $D=0
M1245 168 66 395 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=29630 $D=0
M1246 396 67 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=25000 $D=0
M1247 397 67 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=29630 $D=0
M1248 398 394 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=25000 $D=0
M1249 399 395 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=29630 $D=0
M1250 167 398 735 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=25000 $D=0
M1251 168 399 736 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=29630 $D=0
M1252 400 735 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=25000 $D=0
M1253 401 736 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=29630 $D=0
M1254 398 66 400 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=25000 $D=0
M1255 399 66 401 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=29630 $D=0
M1256 400 396 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=25000 $D=0
M1257 401 397 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=29630 $D=0
M1258 242 402 400 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=25000 $D=0
M1259 243 403 401 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=29630 $D=0
M1260 402 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=25000 $D=0
M1261 403 68 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=29630 $D=0
M1262 167 69 404 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=25000 $D=0
M1263 168 69 405 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=29630 $D=0
M1264 406 70 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=25000 $D=0
M1265 407 70 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=29630 $D=0
M1266 408 404 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=25000 $D=0
M1267 409 405 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=29630 $D=0
M1268 167 408 737 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=25000 $D=0
M1269 168 409 738 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=29630 $D=0
M1270 410 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=25000 $D=0
M1271 411 738 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=29630 $D=0
M1272 408 69 410 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=25000 $D=0
M1273 409 69 411 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=29630 $D=0
M1274 410 406 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=25000 $D=0
M1275 411 407 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=29630 $D=0
M1276 242 412 410 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=25000 $D=0
M1277 243 413 411 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=29630 $D=0
M1278 412 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=25000 $D=0
M1279 413 71 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=29630 $D=0
M1280 167 72 414 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=25000 $D=0
M1281 168 72 415 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=29630 $D=0
M1282 416 73 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=25000 $D=0
M1283 417 73 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=29630 $D=0
M1284 418 414 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=25000 $D=0
M1285 419 415 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=29630 $D=0
M1286 167 418 739 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=25000 $D=0
M1287 168 419 740 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=29630 $D=0
M1288 420 739 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=25000 $D=0
M1289 421 740 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=29630 $D=0
M1290 418 72 420 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=25000 $D=0
M1291 419 72 421 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=29630 $D=0
M1292 420 416 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=25000 $D=0
M1293 421 417 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=29630 $D=0
M1294 242 422 420 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=25000 $D=0
M1295 243 423 421 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=29630 $D=0
M1296 422 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=25000 $D=0
M1297 423 74 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=29630 $D=0
M1298 167 75 424 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=25000 $D=0
M1299 168 75 425 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=29630 $D=0
M1300 426 76 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=25000 $D=0
M1301 427 76 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=29630 $D=0
M1302 428 424 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=25000 $D=0
M1303 429 425 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=29630 $D=0
M1304 167 428 741 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=25000 $D=0
M1305 168 429 742 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=29630 $D=0
M1306 430 741 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=25000 $D=0
M1307 431 742 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=29630 $D=0
M1308 428 75 430 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=25000 $D=0
M1309 429 75 431 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=29630 $D=0
M1310 430 426 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=25000 $D=0
M1311 431 427 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=29630 $D=0
M1312 242 432 430 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=25000 $D=0
M1313 243 433 431 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=29630 $D=0
M1314 432 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=25000 $D=0
M1315 433 77 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=29630 $D=0
M1316 167 78 434 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=25000 $D=0
M1317 168 78 435 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=29630 $D=0
M1318 436 79 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=25000 $D=0
M1319 437 79 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=29630 $D=0
M1320 438 434 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=25000 $D=0
M1321 439 435 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=29630 $D=0
M1322 167 438 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=25000 $D=0
M1323 168 439 744 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=29630 $D=0
M1324 440 743 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=25000 $D=0
M1325 441 744 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=29630 $D=0
M1326 438 78 440 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=25000 $D=0
M1327 439 78 441 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=29630 $D=0
M1328 440 436 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=25000 $D=0
M1329 441 437 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=29630 $D=0
M1330 242 442 440 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=25000 $D=0
M1331 243 443 441 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=29630 $D=0
M1332 442 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=25000 $D=0
M1333 443 80 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=29630 $D=0
M1334 167 81 444 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=25000 $D=0
M1335 168 81 445 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=29630 $D=0
M1336 446 82 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=25000 $D=0
M1337 447 82 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=29630 $D=0
M1338 448 444 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=25000 $D=0
M1339 449 445 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=29630 $D=0
M1340 167 448 745 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=25000 $D=0
M1341 168 449 746 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=29630 $D=0
M1342 450 745 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=25000 $D=0
M1343 451 746 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=29630 $D=0
M1344 448 81 450 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=25000 $D=0
M1345 449 81 451 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=29630 $D=0
M1346 450 446 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=25000 $D=0
M1347 451 447 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=29630 $D=0
M1348 242 452 450 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=25000 $D=0
M1349 243 453 451 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=29630 $D=0
M1350 452 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=25000 $D=0
M1351 453 83 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=29630 $D=0
M1352 167 84 454 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=25000 $D=0
M1353 168 84 455 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=29630 $D=0
M1354 456 85 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=25000 $D=0
M1355 457 85 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=29630 $D=0
M1356 458 454 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=25000 $D=0
M1357 459 455 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=29630 $D=0
M1358 167 458 747 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=25000 $D=0
M1359 168 459 748 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=29630 $D=0
M1360 460 747 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=25000 $D=0
M1361 461 748 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=29630 $D=0
M1362 458 84 460 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=25000 $D=0
M1363 459 84 461 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=29630 $D=0
M1364 460 456 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=25000 $D=0
M1365 461 457 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=29630 $D=0
M1366 242 462 460 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=25000 $D=0
M1367 243 463 461 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=29630 $D=0
M1368 462 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=25000 $D=0
M1369 463 86 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=29630 $D=0
M1370 167 87 464 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=25000 $D=0
M1371 168 87 465 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=29630 $D=0
M1372 466 88 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=25000 $D=0
M1373 467 88 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=29630 $D=0
M1374 468 464 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=25000 $D=0
M1375 469 465 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=29630 $D=0
M1376 167 468 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=25000 $D=0
M1377 168 469 750 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=29630 $D=0
M1378 470 749 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=25000 $D=0
M1379 471 750 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=29630 $D=0
M1380 468 87 470 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=25000 $D=0
M1381 469 87 471 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=29630 $D=0
M1382 470 466 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=25000 $D=0
M1383 471 467 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=29630 $D=0
M1384 242 472 470 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=25000 $D=0
M1385 243 473 471 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=29630 $D=0
M1386 472 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=25000 $D=0
M1387 473 89 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=29630 $D=0
M1388 167 90 474 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=25000 $D=0
M1389 168 90 475 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=29630 $D=0
M1390 476 91 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=25000 $D=0
M1391 477 91 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=29630 $D=0
M1392 478 474 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=25000 $D=0
M1393 479 475 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=29630 $D=0
M1394 167 478 751 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=25000 $D=0
M1395 168 479 752 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=29630 $D=0
M1396 480 751 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=25000 $D=0
M1397 481 752 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=29630 $D=0
M1398 478 90 480 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=25000 $D=0
M1399 479 90 481 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=29630 $D=0
M1400 480 476 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=25000 $D=0
M1401 481 477 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=29630 $D=0
M1402 242 482 480 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=25000 $D=0
M1403 243 483 481 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=29630 $D=0
M1404 482 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=25000 $D=0
M1405 483 92 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=29630 $D=0
M1406 167 93 484 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=25000 $D=0
M1407 168 93 485 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=29630 $D=0
M1408 486 94 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=25000 $D=0
M1409 487 94 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=29630 $D=0
M1410 488 484 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=25000 $D=0
M1411 489 485 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=29630 $D=0
M1412 167 488 753 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=25000 $D=0
M1413 168 489 754 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=29630 $D=0
M1414 490 753 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=25000 $D=0
M1415 491 754 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=29630 $D=0
M1416 488 93 490 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=25000 $D=0
M1417 489 93 491 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=29630 $D=0
M1418 490 486 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=25000 $D=0
M1419 491 487 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=29630 $D=0
M1420 242 492 490 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=25000 $D=0
M1421 243 493 491 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=29630 $D=0
M1422 492 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=25000 $D=0
M1423 493 95 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=29630 $D=0
M1424 167 96 494 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=25000 $D=0
M1425 168 96 495 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=29630 $D=0
M1426 496 97 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=25000 $D=0
M1427 497 97 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=29630 $D=0
M1428 498 494 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=25000 $D=0
M1429 499 495 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=29630 $D=0
M1430 167 498 755 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=25000 $D=0
M1431 168 499 756 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=29630 $D=0
M1432 500 755 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=25000 $D=0
M1433 501 756 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=29630 $D=0
M1434 498 96 500 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=25000 $D=0
M1435 499 96 501 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=29630 $D=0
M1436 500 496 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=25000 $D=0
M1437 501 497 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=29630 $D=0
M1438 242 502 500 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=25000 $D=0
M1439 243 503 501 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=29630 $D=0
M1440 502 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=25000 $D=0
M1441 503 98 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=29630 $D=0
M1442 167 99 504 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=25000 $D=0
M1443 168 99 505 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=29630 $D=0
M1444 506 100 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=25000 $D=0
M1445 507 100 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=29630 $D=0
M1446 508 504 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=25000 $D=0
M1447 509 505 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=29630 $D=0
M1448 167 508 757 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=25000 $D=0
M1449 168 509 758 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=29630 $D=0
M1450 510 757 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=25000 $D=0
M1451 511 758 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=29630 $D=0
M1452 508 99 510 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=25000 $D=0
M1453 509 99 511 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=29630 $D=0
M1454 510 506 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=25000 $D=0
M1455 511 507 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=29630 $D=0
M1456 242 512 510 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=25000 $D=0
M1457 243 513 511 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=29630 $D=0
M1458 512 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=25000 $D=0
M1459 513 101 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=29630 $D=0
M1460 167 102 514 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=25000 $D=0
M1461 168 102 515 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=29630 $D=0
M1462 516 103 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=25000 $D=0
M1463 517 103 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=29630 $D=0
M1464 518 514 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=25000 $D=0
M1465 519 515 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=29630 $D=0
M1466 167 518 759 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=25000 $D=0
M1467 168 519 760 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=29630 $D=0
M1468 520 759 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=25000 $D=0
M1469 521 760 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=29630 $D=0
M1470 518 102 520 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=25000 $D=0
M1471 519 102 521 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=29630 $D=0
M1472 520 516 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=25000 $D=0
M1473 521 517 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=29630 $D=0
M1474 242 522 520 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=25000 $D=0
M1475 243 523 521 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=29630 $D=0
M1476 522 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=25000 $D=0
M1477 523 104 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=29630 $D=0
M1478 167 105 524 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=25000 $D=0
M1479 168 105 525 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=29630 $D=0
M1480 526 106 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=25000 $D=0
M1481 527 106 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=29630 $D=0
M1482 528 524 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=25000 $D=0
M1483 529 525 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=29630 $D=0
M1484 167 528 761 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=25000 $D=0
M1485 168 529 762 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=29630 $D=0
M1486 530 761 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=25000 $D=0
M1487 531 762 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=29630 $D=0
M1488 528 105 530 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=25000 $D=0
M1489 529 105 531 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=29630 $D=0
M1490 530 526 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=25000 $D=0
M1491 531 527 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=29630 $D=0
M1492 242 532 530 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=25000 $D=0
M1493 243 533 531 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=29630 $D=0
M1494 532 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=25000 $D=0
M1495 533 108 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=29630 $D=0
M1496 167 109 534 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=25000 $D=0
M1497 168 109 535 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=29630 $D=0
M1498 536 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=25000 $D=0
M1499 537 110 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=29630 $D=0
M1500 538 534 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=25000 $D=0
M1501 539 535 229 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=29630 $D=0
M1502 167 538 763 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=25000 $D=0
M1503 168 539 764 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=29630 $D=0
M1504 540 763 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=25000 $D=0
M1505 541 764 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=29630 $D=0
M1506 538 109 540 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=25000 $D=0
M1507 539 109 541 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=29630 $D=0
M1508 540 536 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=25000 $D=0
M1509 541 537 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=29630 $D=0
M1510 242 542 540 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=25000 $D=0
M1511 243 543 541 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=29630 $D=0
M1512 542 112 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=25000 $D=0
M1513 543 112 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=29630 $D=0
M1514 167 113 544 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=25000 $D=0
M1515 168 113 545 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=29630 $D=0
M1516 546 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=25000 $D=0
M1517 547 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=29630 $D=0
M1518 6 546 238 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=25000 $D=0
M1519 7 547 239 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=29630 $D=0
M1520 242 544 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=25000 $D=0
M1521 243 545 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=29630 $D=0
M1522 167 550 548 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=25000 $D=0
M1523 168 551 549 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=29630 $D=0
M1524 550 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=25000 $D=0
M1525 551 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=29630 $D=0
M1526 765 238 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=25000 $D=0
M1527 766 239 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=29630 $D=0
M1528 552 550 765 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=25000 $D=0
M1529 553 551 766 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=29630 $D=0
M1530 167 552 554 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=25000 $D=0
M1531 168 553 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=29630 $D=0
M1532 767 554 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=25000 $D=0
M1533 768 555 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=29630 $D=0
M1534 552 548 767 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=25000 $D=0
M1535 553 549 768 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=29630 $D=0
M1536 167 558 556 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=25000 $D=0
M1537 168 559 557 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=29630 $D=0
M1538 558 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=25000 $D=0
M1539 559 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=29630 $D=0
M1540 769 242 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=25000 $D=0
M1541 770 243 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=29630 $D=0
M1542 560 558 769 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=25000 $D=0
M1543 561 559 770 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=29630 $D=0
M1544 167 560 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=25000 $D=0
M1545 168 561 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=29630 $D=0
M1546 771 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=25000 $D=0
M1547 772 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=29630 $D=0
M1548 560 556 771 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=25000 $D=0
M1549 561 557 772 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=29630 $D=0
M1550 562 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=25000 $D=0
M1551 563 120 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=29630 $D=0
M1552 564 120 554 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=25000 $D=0
M1553 565 120 555 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=29630 $D=0
M1554 121 562 564 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=25000 $D=0
M1555 122 563 565 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=29630 $D=0
M1556 566 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=25000 $D=0
M1557 567 123 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=29630 $D=0
M1558 568 123 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=25000 $D=0
M1559 569 123 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=29630 $D=0
M1560 773 566 568 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=25000 $D=0
M1561 774 567 569 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=29630 $D=0
M1562 167 118 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=25000 $D=0
M1563 168 119 774 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=29630 $D=0
M1564 570 124 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=25000 $D=0
M1565 571 124 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=29630 $D=0
M1566 572 124 568 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=25000 $D=0
M1567 573 124 569 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=29630 $D=0
M1568 12 570 572 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=25000 $D=0
M1569 13 571 573 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=29630 $D=0
M1570 576 574 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=25000 $D=0
M1571 577 575 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=29630 $D=0
M1572 167 580 578 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=25000 $D=0
M1573 168 581 579 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=29630 $D=0
M1574 582 564 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=25000 $D=0
M1575 583 565 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=29630 $D=0
M1576 580 564 574 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=25000 $D=0
M1577 581 565 575 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=29630 $D=0
M1578 576 582 580 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=25000 $D=0
M1579 577 583 581 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=29630 $D=0
M1580 584 578 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=25000 $D=0
M1581 585 579 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=29630 $D=0
M1582 125 578 572 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=25000 $D=0
M1583 574 579 573 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=29630 $D=0
M1584 564 584 125 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=25000 $D=0
M1585 565 585 574 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=29630 $D=0
M1586 586 125 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=25000 $D=0
M1587 587 574 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=29630 $D=0
M1588 588 578 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=25000 $D=0
M1589 589 579 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=29630 $D=0
M1590 590 578 586 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=25000 $D=0
M1591 591 579 587 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=29630 $D=0
M1592 572 588 590 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=25000 $D=0
M1593 573 589 591 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=29630 $D=0
M1594 785 564 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=24640 $D=0
M1595 786 565 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=29270 $D=0
M1596 592 572 785 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=24640 $D=0
M1597 593 573 786 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=29270 $D=0
M1598 594 590 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=25000 $D=0
M1599 595 591 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=29630 $D=0
M1600 596 564 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=25000 $D=0
M1601 597 565 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=29630 $D=0
M1602 167 572 596 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=25000 $D=0
M1603 168 573 597 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=29630 $D=0
M1604 598 564 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=25000 $D=0
M1605 599 565 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=29630 $D=0
M1606 167 572 598 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=25000 $D=0
M1607 168 573 599 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=29630 $D=0
M1608 787 564 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=24820 $D=0
M1609 788 565 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=29450 $D=0
M1610 602 572 787 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=24820 $D=0
M1611 603 573 788 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=29450 $D=0
M1612 167 598 602 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=25000 $D=0
M1613 168 599 603 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=29630 $D=0
M1614 604 128 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=25000 $D=0
M1615 605 128 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=29630 $D=0
M1616 606 128 592 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=25000 $D=0
M1617 607 128 593 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=29630 $D=0
M1618 596 604 606 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=25000 $D=0
M1619 597 605 607 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=29630 $D=0
M1620 608 128 594 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=25000 $D=0
M1621 609 128 595 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=29630 $D=0
M1622 602 604 608 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=25000 $D=0
M1623 603 605 609 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=29630 $D=0
M1624 610 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=25000 $D=0
M1625 611 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=29630 $D=0
M1626 612 129 608 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=25000 $D=0
M1627 613 129 609 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=29630 $D=0
M1628 606 610 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=25000 $D=0
M1629 607 611 613 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=29630 $D=0
M1630 14 612 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=25000 $D=0
M1631 15 613 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=29630 $D=0
M1632 614 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=25000 $D=0
M1633 615 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=29630 $D=0
M1634 616 130 131 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=25000 $D=0
M1635 617 130 132 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=29630 $D=0
M1636 133 614 616 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=25000 $D=0
M1637 134 615 617 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=29630 $D=0
M1638 618 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=25000 $D=0
M1639 619 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=29630 $D=0
M1640 620 130 135 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=25000 $D=0
M1641 621 130 136 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=29630 $D=0
M1642 137 618 620 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=25000 $D=0
M1643 138 619 621 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=29630 $D=0
M1644 622 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=25000 $D=0
M1645 623 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=29630 $D=0
M1646 624 130 127 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=25000 $D=0
M1647 625 130 126 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=29630 $D=0
M1648 139 622 624 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=25000 $D=0
M1649 140 623 625 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=29630 $D=0
M1650 626 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=25000 $D=0
M1651 627 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=29630 $D=0
M1652 628 130 142 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=25000 $D=0
M1653 629 130 143 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=29630 $D=0
M1654 144 626 628 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=25000 $D=0
M1655 144 627 629 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=29630 $D=0
M1656 630 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=25000 $D=0
M1657 631 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=29630 $D=0
M1658 632 130 145 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=25000 $D=0
M1659 633 130 146 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=29630 $D=0
M1660 144 630 632 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=25000 $D=0
M1661 144 631 633 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=29630 $D=0
M1662 167 564 775 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=25000 $D=0
M1663 168 565 776 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=29630 $D=0
M1664 134 775 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=25000 $D=0
M1665 131 776 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=29630 $D=0
M1666 634 147 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=25000 $D=0
M1667 635 147 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=29630 $D=0
M1668 148 147 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=25000 $D=0
M1669 149 147 131 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=29630 $D=0
M1670 616 634 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=25000 $D=0
M1671 617 635 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=29630 $D=0
M1672 636 150 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=25000 $D=0
M1673 637 150 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=29630 $D=0
M1674 151 150 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=25000 $D=0
M1675 107 150 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=29630 $D=0
M1676 620 636 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=25000 $D=0
M1677 621 637 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=29630 $D=0
M1678 638 152 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=25000 $D=0
M1679 639 152 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=29630 $D=0
M1680 153 152 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=25000 $D=0
M1681 115 152 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=29630 $D=0
M1682 624 638 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=25000 $D=0
M1683 625 639 115 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=29630 $D=0
M1684 640 154 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=25000 $D=0
M1685 641 154 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=29630 $D=0
M1686 155 154 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=25000 $D=0
M1687 156 154 115 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=29630 $D=0
M1688 628 640 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=25000 $D=0
M1689 629 641 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=29630 $D=0
M1690 642 157 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=25000 $D=0
M1691 643 157 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=29630 $D=0
M1692 214 157 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=25000 $D=0
M1693 215 157 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=29630 $D=0
M1694 632 642 214 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=25000 $D=0
M1695 633 643 215 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=29630 $D=0
M1696 644 158 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=25000 $D=0
M1697 645 158 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=29630 $D=0
M1698 646 158 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=25000 $D=0
M1699 647 158 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=29630 $D=0
M1700 12 644 646 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=25000 $D=0
M1701 13 645 647 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=29630 $D=0
M1702 648 554 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=25000 $D=0
M1703 649 555 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=29630 $D=0
M1704 167 646 648 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=25000 $D=0
M1705 168 647 649 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=29630 $D=0
M1706 789 554 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=24820 $D=0
M1707 790 555 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=29450 $D=0
M1708 652 646 789 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=24820 $D=0
M1709 653 647 790 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=29450 $D=0
M1710 167 648 652 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=25000 $D=0
M1711 168 649 653 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=29630 $D=0
M1712 777 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=25000 $D=0
M1713 778 654 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=29630 $D=0
M1714 167 652 777 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=25000 $D=0
M1715 168 653 778 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=29630 $D=0
M1716 654 777 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=25000 $D=0
M1717 160 778 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=29630 $D=0
M1718 791 554 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=24640 $D=0
M1719 792 555 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=29270 $D=0
M1720 655 657 791 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=24640 $D=0
M1721 656 658 792 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=29270 $D=0
M1722 657 646 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=25000 $D=0
M1723 658 647 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=29630 $D=0
M1724 659 655 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=25000 $D=0
M1725 660 656 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=29630 $D=0
M1726 167 159 659 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=25000 $D=0
M1727 168 654 660 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=29630 $D=0
M1728 662 161 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=25000 $D=0
M1729 663 661 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=29630 $D=0
M1730 661 659 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=25000 $D=0
M1731 162 660 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=29630 $D=0
M1732 167 662 661 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=25000 $D=0
M1733 168 663 162 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=29630 $D=0
M1734 665 664 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=25000 $D=0
M1735 666 163 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=29630 $D=0
M1736 167 669 667 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=25000 $D=0
M1737 168 670 668 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=29630 $D=0
M1738 671 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=25000 $D=0
M1739 672 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=29630 $D=0
M1740 669 121 664 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=25000 $D=0
M1741 670 122 163 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=29630 $D=0
M1742 665 671 669 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=25000 $D=0
M1743 666 672 670 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=29630 $D=0
M1744 673 667 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=25000 $D=0
M1745 674 668 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=29630 $D=0
M1746 164 667 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=25000 $D=0
M1747 664 668 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=29630 $D=0
M1748 121 673 164 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=25000 $D=0
M1749 122 674 664 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=29630 $D=0
M1750 675 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=25000 $D=0
M1751 676 664 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=29630 $D=0
M1752 677 667 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=25000 $D=0
M1753 678 668 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=29630 $D=0
M1754 216 667 675 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=25000 $D=0
M1755 217 668 676 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=29630 $D=0
M1756 6 677 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=25000 $D=0
M1757 7 678 217 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=29630 $D=0
M1758 679 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=25000 $D=0
M1759 680 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=29630 $D=0
M1760 681 165 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=25000 $D=0
M1761 682 165 217 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=29630 $D=0
M1762 14 679 681 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=25000 $D=0
M1763 15 680 682 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=29630 $D=0
M1764 683 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=25000 $D=0
M1765 684 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=29630 $D=0
M1766 166 166 681 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=25000 $D=0
M1767 166 166 682 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=29630 $D=0
M1768 6 683 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=25000 $D=0
M1769 7 684 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=29630 $D=0
M1770 685 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=25000 $D=0
M1771 686 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=29630 $D=0
M1772 167 685 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=25000 $D=0
M1773 168 686 688 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=29630 $D=0
M1774 689 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=25000 $D=0
M1775 690 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=29630 $D=0
M1776 691 687 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=25000 $D=0
M1777 692 688 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=29630 $D=0
M1778 167 691 779 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=25000 $D=0
M1779 168 692 780 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=29630 $D=0
M1780 693 779 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=25000 $D=0
M1781 694 780 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=29630 $D=0
M1782 691 685 693 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=25000 $D=0
M1783 692 686 694 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=29630 $D=0
M1784 695 689 693 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=25000 $D=0
M1785 696 690 694 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=29630 $D=0
M1786 167 699 697 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=25000 $D=0
M1787 168 700 698 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=29630 $D=0
M1788 699 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=25000 $D=0
M1789 700 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=29630 $D=0
M1790 781 695 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=25000 $D=0
M1791 782 696 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=29630 $D=0
M1792 701 699 781 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=25000 $D=0
M1793 702 700 782 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=29630 $D=0
M1794 167 701 121 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=25000 $D=0
M1795 168 702 122 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=29630 $D=0
M1796 783 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=25000 $D=0
M1797 784 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=29630 $D=0
M1798 701 697 783 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=25000 $D=0
M1799 702 698 784 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=29630 $D=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 110 111 112 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168
** N=797 EP=164 IP=1514 FDC=1800
M0 183 1 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=14490 $D=1
M1 184 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=19120 $D=1
M2 185 183 2 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=14490 $D=1
M3 186 184 3 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=19120 $D=1
M4 6 1 185 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=14490 $D=1
M5 7 1 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=19120 $D=1
M6 187 183 4 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=14490 $D=1
M7 188 184 4 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=19120 $D=1
M8 5 1 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=14490 $D=1
M9 5 1 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=19120 $D=1
M10 189 183 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=14490 $D=1
M11 190 184 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=19120 $D=1
M12 6 1 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=14490 $D=1
M13 7 1 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=19120 $D=1
M14 193 191 189 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=14490 $D=1
M15 194 192 190 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=19120 $D=1
M16 191 9 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=14490 $D=1
M17 192 9 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=19120 $D=1
M18 195 191 187 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=14490 $D=1
M19 196 192 188 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=19120 $D=1
M20 185 9 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=14490 $D=1
M21 186 9 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=19120 $D=1
M22 197 10 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=14490 $D=1
M23 198 10 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=19120 $D=1
M24 199 197 195 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=14490 $D=1
M25 200 198 196 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=19120 $D=1
M26 193 10 199 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=14490 $D=1
M27 194 10 200 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=19120 $D=1
M28 201 11 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=14490 $D=1
M29 202 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=19120 $D=1
M30 203 201 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=14490 $D=1
M31 204 202 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=19120 $D=1
M32 12 11 203 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=14490 $D=1
M33 13 11 204 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=19120 $D=1
M34 205 201 14 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=14490 $D=1
M35 206 202 15 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=19120 $D=1
M36 207 11 205 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=14490 $D=1
M37 208 11 206 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=19120 $D=1
M38 211 201 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=14490 $D=1
M39 212 202 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=19120 $D=1
M40 199 11 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=14490 $D=1
M41 200 11 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=19120 $D=1
M42 215 213 211 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=14490 $D=1
M43 216 214 212 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=19120 $D=1
M44 213 16 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=14490 $D=1
M45 214 16 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=19120 $D=1
M46 217 213 205 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=14490 $D=1
M47 218 214 206 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=19120 $D=1
M48 203 16 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=14490 $D=1
M49 204 16 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=19120 $D=1
M50 219 17 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=14490 $D=1
M51 220 17 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=19120 $D=1
M52 221 219 217 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=14490 $D=1
M53 222 220 218 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=19120 $D=1
M54 215 17 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=14490 $D=1
M55 216 17 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=19120 $D=1
M56 6 18 223 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=14490 $D=1
M57 7 18 224 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=19120 $D=1
M58 225 19 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=14490 $D=1
M59 226 19 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=19120 $D=1
M60 227 18 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=14490 $D=1
M61 228 18 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=19120 $D=1
M62 6 227 696 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=14490 $D=1
M63 7 228 697 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=19120 $D=1
M64 229 696 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=14490 $D=1
M65 230 697 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=19120 $D=1
M66 227 223 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=14490 $D=1
M67 228 224 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=19120 $D=1
M68 229 19 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=14490 $D=1
M69 230 19 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=19120 $D=1
M70 235 20 229 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=14490 $D=1
M71 236 20 230 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=19120 $D=1
M72 233 20 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=14490 $D=1
M73 234 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=19120 $D=1
M74 6 21 237 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=14490 $D=1
M75 7 21 238 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=19120 $D=1
M76 239 22 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=14490 $D=1
M77 240 22 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=19120 $D=1
M78 241 21 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=14490 $D=1
M79 242 21 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=19120 $D=1
M80 6 241 698 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=14490 $D=1
M81 7 242 699 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=19120 $D=1
M82 243 698 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=14490 $D=1
M83 244 699 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=19120 $D=1
M84 241 237 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=14490 $D=1
M85 242 238 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=19120 $D=1
M86 243 22 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=14490 $D=1
M87 244 22 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=19120 $D=1
M88 235 23 243 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=14490 $D=1
M89 236 23 244 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=19120 $D=1
M90 245 23 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=14490 $D=1
M91 246 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=19120 $D=1
M92 6 24 247 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=14490 $D=1
M93 7 24 248 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=19120 $D=1
M94 249 25 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=14490 $D=1
M95 250 25 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=19120 $D=1
M96 251 24 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=14490 $D=1
M97 252 24 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=19120 $D=1
M98 6 251 700 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=14490 $D=1
M99 7 252 701 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=19120 $D=1
M100 253 700 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=14490 $D=1
M101 254 701 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=19120 $D=1
M102 251 247 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=14490 $D=1
M103 252 248 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=19120 $D=1
M104 253 25 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=14490 $D=1
M105 254 25 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=19120 $D=1
M106 235 26 253 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=14490 $D=1
M107 236 26 254 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=19120 $D=1
M108 255 26 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=14490 $D=1
M109 256 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=19120 $D=1
M110 6 27 257 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=14490 $D=1
M111 7 27 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=19120 $D=1
M112 259 28 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=14490 $D=1
M113 260 28 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=19120 $D=1
M114 261 27 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=14490 $D=1
M115 262 27 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=19120 $D=1
M116 6 261 702 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=14490 $D=1
M117 7 262 703 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=19120 $D=1
M118 263 702 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=14490 $D=1
M119 264 703 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=19120 $D=1
M120 261 257 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=14490 $D=1
M121 262 258 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=19120 $D=1
M122 263 28 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=14490 $D=1
M123 264 28 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=19120 $D=1
M124 235 29 263 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=14490 $D=1
M125 236 29 264 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=19120 $D=1
M126 265 29 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=14490 $D=1
M127 266 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=19120 $D=1
M128 6 30 267 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=14490 $D=1
M129 7 30 268 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=19120 $D=1
M130 269 31 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=14490 $D=1
M131 270 31 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=19120 $D=1
M132 271 30 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=14490 $D=1
M133 272 30 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=19120 $D=1
M134 6 271 704 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=14490 $D=1
M135 7 272 705 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=19120 $D=1
M136 273 704 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=14490 $D=1
M137 274 705 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=19120 $D=1
M138 271 267 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=14490 $D=1
M139 272 268 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=19120 $D=1
M140 273 31 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=14490 $D=1
M141 274 31 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=19120 $D=1
M142 235 32 273 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=14490 $D=1
M143 236 32 274 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=19120 $D=1
M144 275 32 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=14490 $D=1
M145 276 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=19120 $D=1
M146 6 33 277 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=14490 $D=1
M147 7 33 278 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=19120 $D=1
M148 279 34 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=14490 $D=1
M149 280 34 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=19120 $D=1
M150 281 33 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=14490 $D=1
M151 282 33 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=19120 $D=1
M152 6 281 706 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=14490 $D=1
M153 7 282 707 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=19120 $D=1
M154 283 706 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=14490 $D=1
M155 284 707 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=19120 $D=1
M156 281 277 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=14490 $D=1
M157 282 278 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=19120 $D=1
M158 283 34 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=14490 $D=1
M159 284 34 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=19120 $D=1
M160 235 35 283 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=14490 $D=1
M161 236 35 284 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=19120 $D=1
M162 285 35 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=14490 $D=1
M163 286 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=19120 $D=1
M164 6 36 287 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=14490 $D=1
M165 7 36 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=19120 $D=1
M166 289 37 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=14490 $D=1
M167 290 37 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=19120 $D=1
M168 291 36 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=14490 $D=1
M169 292 36 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=19120 $D=1
M170 6 291 708 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=14490 $D=1
M171 7 292 709 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=19120 $D=1
M172 293 708 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=14490 $D=1
M173 294 709 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=19120 $D=1
M174 291 287 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=14490 $D=1
M175 292 288 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=19120 $D=1
M176 293 37 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=14490 $D=1
M177 294 37 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=19120 $D=1
M178 235 38 293 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=14490 $D=1
M179 236 38 294 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=19120 $D=1
M180 295 38 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=14490 $D=1
M181 296 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=19120 $D=1
M182 6 39 297 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=14490 $D=1
M183 7 39 298 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=19120 $D=1
M184 299 40 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=14490 $D=1
M185 300 40 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=19120 $D=1
M186 301 39 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=14490 $D=1
M187 302 39 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=19120 $D=1
M188 6 301 710 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=14490 $D=1
M189 7 302 711 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=19120 $D=1
M190 303 710 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=14490 $D=1
M191 304 711 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=19120 $D=1
M192 301 297 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=14490 $D=1
M193 302 298 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=19120 $D=1
M194 303 40 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=14490 $D=1
M195 304 40 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=19120 $D=1
M196 235 41 303 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=14490 $D=1
M197 236 41 304 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=19120 $D=1
M198 305 41 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=14490 $D=1
M199 306 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=19120 $D=1
M200 6 42 307 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=14490 $D=1
M201 7 42 308 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=19120 $D=1
M202 309 43 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=14490 $D=1
M203 310 43 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=19120 $D=1
M204 311 42 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=14490 $D=1
M205 312 42 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=19120 $D=1
M206 6 311 712 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=14490 $D=1
M207 7 312 713 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=19120 $D=1
M208 313 712 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=14490 $D=1
M209 314 713 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=19120 $D=1
M210 311 307 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=14490 $D=1
M211 312 308 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=19120 $D=1
M212 313 43 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=14490 $D=1
M213 314 43 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=19120 $D=1
M214 235 44 313 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=14490 $D=1
M215 236 44 314 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=19120 $D=1
M216 315 44 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=14490 $D=1
M217 316 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=19120 $D=1
M218 6 45 317 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=14490 $D=1
M219 7 45 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=19120 $D=1
M220 319 46 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=14490 $D=1
M221 320 46 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=19120 $D=1
M222 321 45 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=14490 $D=1
M223 322 45 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=19120 $D=1
M224 6 321 714 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=14490 $D=1
M225 7 322 715 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=19120 $D=1
M226 323 714 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=14490 $D=1
M227 324 715 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=19120 $D=1
M228 321 317 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=14490 $D=1
M229 322 318 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=19120 $D=1
M230 323 46 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=14490 $D=1
M231 324 46 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=19120 $D=1
M232 235 47 323 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=14490 $D=1
M233 236 47 324 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=19120 $D=1
M234 325 47 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=14490 $D=1
M235 326 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=19120 $D=1
M236 6 48 327 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=14490 $D=1
M237 7 48 328 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=19120 $D=1
M238 329 49 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=14490 $D=1
M239 330 49 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=19120 $D=1
M240 331 48 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=14490 $D=1
M241 332 48 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=19120 $D=1
M242 6 331 716 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=14490 $D=1
M243 7 332 717 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=19120 $D=1
M244 333 716 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=14490 $D=1
M245 334 717 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=19120 $D=1
M246 331 327 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=14490 $D=1
M247 332 328 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=19120 $D=1
M248 333 49 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=14490 $D=1
M249 334 49 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=19120 $D=1
M250 235 50 333 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=14490 $D=1
M251 236 50 334 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=19120 $D=1
M252 335 50 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=14490 $D=1
M253 336 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=19120 $D=1
M254 6 51 337 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=14490 $D=1
M255 7 51 338 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=19120 $D=1
M256 339 52 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=14490 $D=1
M257 340 52 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=19120 $D=1
M258 341 51 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=14490 $D=1
M259 342 51 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=19120 $D=1
M260 6 341 718 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=14490 $D=1
M261 7 342 719 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=19120 $D=1
M262 343 718 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=14490 $D=1
M263 344 719 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=19120 $D=1
M264 341 337 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=14490 $D=1
M265 342 338 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=19120 $D=1
M266 343 52 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=14490 $D=1
M267 344 52 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=19120 $D=1
M268 235 53 343 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=14490 $D=1
M269 236 53 344 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=19120 $D=1
M270 345 53 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=14490 $D=1
M271 346 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=19120 $D=1
M272 6 54 347 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=14490 $D=1
M273 7 54 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=19120 $D=1
M274 349 55 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=14490 $D=1
M275 350 55 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=19120 $D=1
M276 351 54 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=14490 $D=1
M277 352 54 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=19120 $D=1
M278 6 351 720 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=14490 $D=1
M279 7 352 721 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=19120 $D=1
M280 353 720 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=14490 $D=1
M281 354 721 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=19120 $D=1
M282 351 347 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=14490 $D=1
M283 352 348 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=19120 $D=1
M284 353 55 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=14490 $D=1
M285 354 55 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=19120 $D=1
M286 235 56 353 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=14490 $D=1
M287 236 56 354 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=19120 $D=1
M288 355 56 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=14490 $D=1
M289 356 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=19120 $D=1
M290 6 57 357 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=14490 $D=1
M291 7 57 358 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=19120 $D=1
M292 359 58 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=14490 $D=1
M293 360 58 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=19120 $D=1
M294 361 57 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=14490 $D=1
M295 362 57 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=19120 $D=1
M296 6 361 722 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=14490 $D=1
M297 7 362 723 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=19120 $D=1
M298 363 722 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=14490 $D=1
M299 364 723 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=19120 $D=1
M300 361 357 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=14490 $D=1
M301 362 358 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=19120 $D=1
M302 363 58 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=14490 $D=1
M303 364 58 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=19120 $D=1
M304 235 59 363 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=14490 $D=1
M305 236 59 364 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=19120 $D=1
M306 365 59 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=14490 $D=1
M307 366 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=19120 $D=1
M308 6 60 367 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=14490 $D=1
M309 7 60 368 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=19120 $D=1
M310 369 61 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=14490 $D=1
M311 370 61 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=19120 $D=1
M312 371 60 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=14490 $D=1
M313 372 60 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=19120 $D=1
M314 6 371 724 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=14490 $D=1
M315 7 372 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=19120 $D=1
M316 373 724 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=14490 $D=1
M317 374 725 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=19120 $D=1
M318 371 367 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=14490 $D=1
M319 372 368 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=19120 $D=1
M320 373 61 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=14490 $D=1
M321 374 61 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=19120 $D=1
M322 235 62 373 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=14490 $D=1
M323 236 62 374 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=19120 $D=1
M324 375 62 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=14490 $D=1
M325 376 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=19120 $D=1
M326 6 63 377 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=14490 $D=1
M327 7 63 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=19120 $D=1
M328 379 64 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=14490 $D=1
M329 380 64 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=19120 $D=1
M330 381 63 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=14490 $D=1
M331 382 63 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=19120 $D=1
M332 6 381 726 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=14490 $D=1
M333 7 382 727 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=19120 $D=1
M334 383 726 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=14490 $D=1
M335 384 727 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=19120 $D=1
M336 381 377 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=14490 $D=1
M337 382 378 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=19120 $D=1
M338 383 64 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=14490 $D=1
M339 384 64 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=19120 $D=1
M340 235 65 383 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=14490 $D=1
M341 236 65 384 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=19120 $D=1
M342 385 65 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=14490 $D=1
M343 386 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=19120 $D=1
M344 6 66 387 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=14490 $D=1
M345 7 66 388 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=19120 $D=1
M346 389 67 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=14490 $D=1
M347 390 67 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=19120 $D=1
M348 391 66 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=14490 $D=1
M349 392 66 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=19120 $D=1
M350 6 391 728 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=14490 $D=1
M351 7 392 729 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=19120 $D=1
M352 393 728 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=14490 $D=1
M353 394 729 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=19120 $D=1
M354 391 387 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=14490 $D=1
M355 392 388 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=19120 $D=1
M356 393 67 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=14490 $D=1
M357 394 67 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=19120 $D=1
M358 235 68 393 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=14490 $D=1
M359 236 68 394 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=19120 $D=1
M360 395 68 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=14490 $D=1
M361 396 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=19120 $D=1
M362 6 69 397 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=14490 $D=1
M363 7 69 398 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=19120 $D=1
M364 399 70 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=14490 $D=1
M365 400 70 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=19120 $D=1
M366 401 69 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=14490 $D=1
M367 402 69 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=19120 $D=1
M368 6 401 730 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=14490 $D=1
M369 7 402 731 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=19120 $D=1
M370 403 730 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=14490 $D=1
M371 404 731 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=19120 $D=1
M372 401 397 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=14490 $D=1
M373 402 398 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=19120 $D=1
M374 403 70 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=14490 $D=1
M375 404 70 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=19120 $D=1
M376 235 71 403 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=14490 $D=1
M377 236 71 404 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=19120 $D=1
M378 405 71 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=14490 $D=1
M379 406 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=19120 $D=1
M380 6 72 407 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=14490 $D=1
M381 7 72 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=19120 $D=1
M382 409 73 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=14490 $D=1
M383 410 73 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=19120 $D=1
M384 411 72 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=14490 $D=1
M385 412 72 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=19120 $D=1
M386 6 411 732 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=14490 $D=1
M387 7 412 733 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=19120 $D=1
M388 413 732 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=14490 $D=1
M389 414 733 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=19120 $D=1
M390 411 407 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=14490 $D=1
M391 412 408 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=19120 $D=1
M392 413 73 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=14490 $D=1
M393 414 73 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=19120 $D=1
M394 235 74 413 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=14490 $D=1
M395 236 74 414 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=19120 $D=1
M396 415 74 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=14490 $D=1
M397 416 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=19120 $D=1
M398 6 75 417 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=14490 $D=1
M399 7 75 418 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=19120 $D=1
M400 419 76 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=14490 $D=1
M401 420 76 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=19120 $D=1
M402 421 75 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=14490 $D=1
M403 422 75 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=19120 $D=1
M404 6 421 734 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=14490 $D=1
M405 7 422 735 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=19120 $D=1
M406 423 734 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=14490 $D=1
M407 424 735 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=19120 $D=1
M408 421 417 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=14490 $D=1
M409 422 418 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=19120 $D=1
M410 423 76 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=14490 $D=1
M411 424 76 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=19120 $D=1
M412 235 77 423 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=14490 $D=1
M413 236 77 424 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=19120 $D=1
M414 425 77 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=14490 $D=1
M415 426 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=19120 $D=1
M416 6 78 427 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=14490 $D=1
M417 7 78 428 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=19120 $D=1
M418 429 79 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=14490 $D=1
M419 430 79 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=19120 $D=1
M420 431 78 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=14490 $D=1
M421 432 78 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=19120 $D=1
M422 6 431 736 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=14490 $D=1
M423 7 432 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=19120 $D=1
M424 433 736 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=14490 $D=1
M425 434 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=19120 $D=1
M426 431 427 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=14490 $D=1
M427 432 428 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=19120 $D=1
M428 433 79 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=14490 $D=1
M429 434 79 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=19120 $D=1
M430 235 80 433 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=14490 $D=1
M431 236 80 434 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=19120 $D=1
M432 435 80 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=14490 $D=1
M433 436 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=19120 $D=1
M434 6 81 437 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=14490 $D=1
M435 7 81 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=19120 $D=1
M436 439 82 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=14490 $D=1
M437 440 82 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=19120 $D=1
M438 441 81 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=14490 $D=1
M439 442 81 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=19120 $D=1
M440 6 441 738 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=14490 $D=1
M441 7 442 739 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=19120 $D=1
M442 443 738 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=14490 $D=1
M443 444 739 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=19120 $D=1
M444 441 437 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=14490 $D=1
M445 442 438 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=19120 $D=1
M446 443 82 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=14490 $D=1
M447 444 82 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=19120 $D=1
M448 235 83 443 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=14490 $D=1
M449 236 83 444 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=19120 $D=1
M450 445 83 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=14490 $D=1
M451 446 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=19120 $D=1
M452 6 84 447 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=14490 $D=1
M453 7 84 448 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=19120 $D=1
M454 449 85 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=14490 $D=1
M455 450 85 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=19120 $D=1
M456 451 84 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=14490 $D=1
M457 452 84 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=19120 $D=1
M458 6 451 740 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=14490 $D=1
M459 7 452 741 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=19120 $D=1
M460 453 740 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=14490 $D=1
M461 454 741 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=19120 $D=1
M462 451 447 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=14490 $D=1
M463 452 448 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=19120 $D=1
M464 453 85 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=14490 $D=1
M465 454 85 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=19120 $D=1
M466 235 86 453 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=14490 $D=1
M467 236 86 454 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=19120 $D=1
M468 455 86 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=14490 $D=1
M469 456 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=19120 $D=1
M470 6 87 457 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=14490 $D=1
M471 7 87 458 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=19120 $D=1
M472 459 88 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=14490 $D=1
M473 460 88 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=19120 $D=1
M474 461 87 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=14490 $D=1
M475 462 87 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=19120 $D=1
M476 6 461 742 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=14490 $D=1
M477 7 462 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=19120 $D=1
M478 463 742 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=14490 $D=1
M479 464 743 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=19120 $D=1
M480 461 457 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=14490 $D=1
M481 462 458 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=19120 $D=1
M482 463 88 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=14490 $D=1
M483 464 88 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=19120 $D=1
M484 235 89 463 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=14490 $D=1
M485 236 89 464 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=19120 $D=1
M486 465 89 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=14490 $D=1
M487 466 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=19120 $D=1
M488 6 90 467 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=14490 $D=1
M489 7 90 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=19120 $D=1
M490 469 91 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=14490 $D=1
M491 470 91 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=19120 $D=1
M492 471 90 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=14490 $D=1
M493 472 90 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=19120 $D=1
M494 6 471 744 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=14490 $D=1
M495 7 472 745 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=19120 $D=1
M496 473 744 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=14490 $D=1
M497 474 745 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=19120 $D=1
M498 471 467 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=14490 $D=1
M499 472 468 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=19120 $D=1
M500 473 91 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=14490 $D=1
M501 474 91 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=19120 $D=1
M502 235 92 473 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=14490 $D=1
M503 236 92 474 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=19120 $D=1
M504 475 92 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=14490 $D=1
M505 476 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=19120 $D=1
M506 6 93 477 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=14490 $D=1
M507 7 93 478 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=19120 $D=1
M508 479 94 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=14490 $D=1
M509 480 94 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=19120 $D=1
M510 481 93 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=14490 $D=1
M511 482 93 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=19120 $D=1
M512 6 481 746 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=14490 $D=1
M513 7 482 747 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=19120 $D=1
M514 483 746 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=14490 $D=1
M515 484 747 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=19120 $D=1
M516 481 477 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=14490 $D=1
M517 482 478 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=19120 $D=1
M518 483 94 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=14490 $D=1
M519 484 94 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=19120 $D=1
M520 235 95 483 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=14490 $D=1
M521 236 95 484 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=19120 $D=1
M522 485 95 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=14490 $D=1
M523 486 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=19120 $D=1
M524 6 96 487 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=14490 $D=1
M525 7 96 488 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=19120 $D=1
M526 489 97 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=14490 $D=1
M527 490 97 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=19120 $D=1
M528 491 96 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=14490 $D=1
M529 492 96 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=19120 $D=1
M530 6 491 748 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=14490 $D=1
M531 7 492 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=19120 $D=1
M532 493 748 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=14490 $D=1
M533 494 749 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=19120 $D=1
M534 491 487 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=14490 $D=1
M535 492 488 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=19120 $D=1
M536 493 97 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=14490 $D=1
M537 494 97 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=19120 $D=1
M538 235 98 493 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=14490 $D=1
M539 236 98 494 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=19120 $D=1
M540 495 98 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=14490 $D=1
M541 496 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=19120 $D=1
M542 6 99 497 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=14490 $D=1
M543 7 99 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=19120 $D=1
M544 499 100 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=14490 $D=1
M545 500 100 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=19120 $D=1
M546 501 99 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=14490 $D=1
M547 502 99 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=19120 $D=1
M548 6 501 750 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=14490 $D=1
M549 7 502 751 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=19120 $D=1
M550 503 750 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=14490 $D=1
M551 504 751 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=19120 $D=1
M552 501 497 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=14490 $D=1
M553 502 498 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=19120 $D=1
M554 503 100 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=14490 $D=1
M555 504 100 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=19120 $D=1
M556 235 101 503 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=14490 $D=1
M557 236 101 504 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=19120 $D=1
M558 505 101 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=14490 $D=1
M559 506 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=19120 $D=1
M560 6 102 507 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=14490 $D=1
M561 7 102 508 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=19120 $D=1
M562 509 103 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=14490 $D=1
M563 510 103 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=19120 $D=1
M564 511 102 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=14490 $D=1
M565 512 102 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=19120 $D=1
M566 6 511 752 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=14490 $D=1
M567 7 512 753 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=19120 $D=1
M568 513 752 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=14490 $D=1
M569 514 753 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=19120 $D=1
M570 511 507 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=14490 $D=1
M571 512 508 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=19120 $D=1
M572 513 103 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=14490 $D=1
M573 514 103 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=19120 $D=1
M574 235 104 513 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=14490 $D=1
M575 236 104 514 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=19120 $D=1
M576 515 104 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=14490 $D=1
M577 516 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=19120 $D=1
M578 6 105 517 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=14490 $D=1
M579 7 105 518 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=19120 $D=1
M580 519 106 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=14490 $D=1
M581 520 106 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=19120 $D=1
M582 521 105 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=14490 $D=1
M583 522 105 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=19120 $D=1
M584 6 521 754 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=14490 $D=1
M585 7 522 755 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=19120 $D=1
M586 523 754 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=14490 $D=1
M587 524 755 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=19120 $D=1
M588 521 517 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=14490 $D=1
M589 522 518 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=19120 $D=1
M590 523 106 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=14490 $D=1
M591 524 106 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=19120 $D=1
M592 235 108 523 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=14490 $D=1
M593 236 108 524 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=19120 $D=1
M594 525 108 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=14490 $D=1
M595 526 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=19120 $D=1
M596 6 110 527 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=14490 $D=1
M597 7 110 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=19120 $D=1
M598 529 111 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=14490 $D=1
M599 530 111 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=19120 $D=1
M600 531 110 221 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=14490 $D=1
M601 532 110 222 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=19120 $D=1
M602 6 531 756 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=14490 $D=1
M603 7 532 757 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=19120 $D=1
M604 533 756 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=14490 $D=1
M605 534 757 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=19120 $D=1
M606 531 527 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=14490 $D=1
M607 532 528 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=19120 $D=1
M608 533 111 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=14490 $D=1
M609 534 111 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=19120 $D=1
M610 235 114 533 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=14490 $D=1
M611 236 114 534 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=19120 $D=1
M612 535 114 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=14490 $D=1
M613 536 114 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=19120 $D=1
M614 6 115 537 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=14490 $D=1
M615 7 115 538 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=19120 $D=1
M616 539 116 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=14490 $D=1
M617 540 116 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=19120 $D=1
M618 6 116 231 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=14490 $D=1
M619 7 116 232 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=19120 $D=1
M620 235 115 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=14490 $D=1
M621 236 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=19120 $D=1
M622 6 543 541 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=14490 $D=1
M623 7 544 542 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=19120 $D=1
M624 543 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=14490 $D=1
M625 544 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=19120 $D=1
M626 758 231 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=14490 $D=1
M627 759 232 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=19120 $D=1
M628 545 541 758 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=14490 $D=1
M629 546 542 759 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=19120 $D=1
M630 6 545 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=14490 $D=1
M631 7 546 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=19120 $D=1
M632 760 547 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=14490 $D=1
M633 761 548 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=19120 $D=1
M634 545 543 760 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=14490 $D=1
M635 546 544 761 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=19120 $D=1
M636 6 551 549 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=14490 $D=1
M637 7 552 550 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=19120 $D=1
M638 551 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=14490 $D=1
M639 552 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=19120 $D=1
M640 762 235 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=14490 $D=1
M641 763 236 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=19120 $D=1
M642 553 549 762 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=14490 $D=1
M643 554 550 763 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=19120 $D=1
M644 6 553 118 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=14490 $D=1
M645 7 554 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=19120 $D=1
M646 764 118 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=14490 $D=1
M647 765 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=19120 $D=1
M648 553 551 764 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=14490 $D=1
M649 554 552 765 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=19120 $D=1
M650 555 120 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=14490 $D=1
M651 556 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=19120 $D=1
M652 557 555 547 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=14490 $D=1
M653 558 556 548 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=19120 $D=1
M654 121 120 557 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=14490 $D=1
M655 122 120 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=19120 $D=1
M656 559 123 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=14490 $D=1
M657 560 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=19120 $D=1
M658 562 559 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=14490 $D=1
M659 563 560 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=19120 $D=1
M660 766 123 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=14490 $D=1
M661 767 123 563 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=19120 $D=1
M662 6 561 766 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=14490 $D=1
M663 7 119 767 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=19120 $D=1
M664 564 124 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=14490 $D=1
M665 565 124 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=19120 $D=1
M666 566 564 562 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=14490 $D=1
M667 567 565 563 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=19120 $D=1
M668 12 124 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=14490 $D=1
M669 13 124 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=19120 $D=1
M670 569 568 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=14490 $D=1
M671 570 125 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=19120 $D=1
M672 6 573 571 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=14490 $D=1
M673 7 574 572 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=19120 $D=1
M674 575 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=14490 $D=1
M675 576 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=19120 $D=1
M676 573 575 568 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=14490 $D=1
M677 574 576 125 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=19120 $D=1
M678 569 557 573 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=14490 $D=1
M679 570 558 574 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=19120 $D=1
M680 577 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=14490 $D=1
M681 578 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=19120 $D=1
M682 126 577 566 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=14490 $D=1
M683 568 578 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=19120 $D=1
M684 557 571 126 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=14490 $D=1
M685 558 572 568 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=19120 $D=1
M686 579 126 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=14490 $D=1
M687 580 568 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=19120 $D=1
M688 581 571 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=14490 $D=1
M689 582 572 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=19120 $D=1
M690 583 581 579 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=14490 $D=1
M691 584 582 580 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=19120 $D=1
M692 566 571 583 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=14490 $D=1
M693 567 572 584 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=19120 $D=1
M694 585 557 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=14490 $D=1
M695 586 558 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=19120 $D=1
M696 6 566 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=14490 $D=1
M697 7 567 586 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=19120 $D=1
M698 587 583 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=14490 $D=1
M699 588 584 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=19120 $D=1
M700 786 557 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=14490 $D=1
M701 787 558 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=19120 $D=1
M702 589 566 786 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=14490 $D=1
M703 590 567 787 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=19120 $D=1
M704 788 557 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=14490 $D=1
M705 789 558 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=19120 $D=1
M706 591 566 788 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=14490 $D=1
M707 592 567 789 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=19120 $D=1
M708 595 557 593 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=14490 $D=1
M709 596 558 594 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=19120 $D=1
M710 593 566 595 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=14490 $D=1
M711 594 567 596 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=19120 $D=1
M712 6 591 593 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=14490 $D=1
M713 7 592 594 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=19120 $D=1
M714 597 129 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=14490 $D=1
M715 598 129 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=19120 $D=1
M716 599 597 585 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=14490 $D=1
M717 600 598 586 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=19120 $D=1
M718 589 129 599 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=14490 $D=1
M719 590 129 600 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=19120 $D=1
M720 601 597 587 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=14490 $D=1
M721 602 598 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=19120 $D=1
M722 595 129 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=14490 $D=1
M723 596 129 602 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=19120 $D=1
M724 603 130 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=14490 $D=1
M725 604 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=19120 $D=1
M726 605 603 601 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=14490 $D=1
M727 606 604 602 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=19120 $D=1
M728 599 130 605 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=14490 $D=1
M729 600 130 606 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=19120 $D=1
M730 14 605 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=14490 $D=1
M731 15 606 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=19120 $D=1
M732 607 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=14490 $D=1
M733 608 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=19120 $D=1
M734 609 607 132 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=14490 $D=1
M735 610 608 133 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=19120 $D=1
M736 134 131 609 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=14490 $D=1
M737 135 131 610 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=19120 $D=1
M738 611 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=14490 $D=1
M739 612 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=19120 $D=1
M740 613 611 136 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=14490 $D=1
M741 614 612 137 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=19120 $D=1
M742 138 131 613 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=14490 $D=1
M743 139 131 614 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=19120 $D=1
M744 615 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=14490 $D=1
M745 616 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=19120 $D=1
M746 617 615 127 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=14490 $D=1
M747 618 616 128 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=19120 $D=1
M748 140 131 617 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=14490 $D=1
M749 141 131 618 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=19120 $D=1
M750 619 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=14490 $D=1
M751 620 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=19120 $D=1
M752 621 619 143 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=14490 $D=1
M753 622 620 144 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=19120 $D=1
M754 140 131 621 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=14490 $D=1
M755 140 131 622 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=19120 $D=1
M756 623 131 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=14490 $D=1
M757 624 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=19120 $D=1
M758 625 623 145 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=14490 $D=1
M759 626 624 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=19120 $D=1
M760 140 131 625 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=14490 $D=1
M761 140 131 626 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=19120 $D=1
M762 6 557 768 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=14490 $D=1
M763 7 558 769 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=19120 $D=1
M764 135 768 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=14490 $D=1
M765 132 769 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=19120 $D=1
M766 627 147 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=14490 $D=1
M767 628 147 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=19120 $D=1
M768 148 627 135 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=14490 $D=1
M769 149 628 132 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=19120 $D=1
M770 609 147 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=14490 $D=1
M771 610 147 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=19120 $D=1
M772 629 150 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=14490 $D=1
M773 630 150 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=19120 $D=1
M774 151 629 148 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=14490 $D=1
M775 107 630 149 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=19120 $D=1
M776 613 150 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=14490 $D=1
M777 614 150 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=19120 $D=1
M778 631 152 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=14490 $D=1
M779 632 152 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=19120 $D=1
M780 153 631 151 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=14490 $D=1
M781 112 632 107 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=19120 $D=1
M782 617 152 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=14490 $D=1
M783 618 152 112 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=19120 $D=1
M784 633 154 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=14490 $D=1
M785 634 154 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=19120 $D=1
M786 155 633 153 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=14490 $D=1
M787 156 634 112 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=19120 $D=1
M788 621 154 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=14490 $D=1
M789 622 154 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=19120 $D=1
M790 635 157 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=14490 $D=1
M791 636 157 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=19120 $D=1
M792 207 635 155 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=14490 $D=1
M793 208 636 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=19120 $D=1
M794 625 157 207 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=14490 $D=1
M795 626 157 208 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=19120 $D=1
M796 637 158 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=14490 $D=1
M797 638 158 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=19120 $D=1
M798 639 637 561 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=14490 $D=1
M799 640 638 119 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=19120 $D=1
M800 12 158 639 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=14490 $D=1
M801 13 158 640 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=19120 $D=1
M802 790 547 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=14490 $D=1
M803 791 548 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=19120 $D=1
M804 641 639 790 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=14490 $D=1
M805 642 640 791 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=19120 $D=1
M806 645 547 643 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=14490 $D=1
M807 646 548 644 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=19120 $D=1
M808 643 639 645 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=14490 $D=1
M809 644 640 646 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=19120 $D=1
M810 6 641 643 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=14490 $D=1
M811 7 642 644 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=19120 $D=1
M812 792 159 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=14490 $D=1
M813 793 647 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=19120 $D=1
M814 770 645 792 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=14490 $D=1
M815 771 646 793 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=19120 $D=1
M816 647 770 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=14490 $D=1
M817 160 771 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=19120 $D=1
M818 648 547 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=14490 $D=1
M819 649 548 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=19120 $D=1
M820 6 650 648 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=14490 $D=1
M821 7 651 649 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=19120 $D=1
M822 650 639 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=14490 $D=1
M823 651 640 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=19120 $D=1
M824 794 648 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=14490 $D=1
M825 795 649 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=19120 $D=1
M826 652 159 794 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=14490 $D=1
M827 653 647 795 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=19120 $D=1
M828 655 161 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=14490 $D=1
M829 656 654 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=19120 $D=1
M830 796 652 6 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=14490 $D=1
M831 797 653 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=19120 $D=1
M832 654 655 796 6 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=14490 $D=1
M833 162 656 797 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=19120 $D=1
M834 658 657 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=14490 $D=1
M835 659 163 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=19120 $D=1
M836 6 662 660 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=14490 $D=1
M837 7 663 661 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=19120 $D=1
M838 664 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=14490 $D=1
M839 665 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=19120 $D=1
M840 662 664 657 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=14490 $D=1
M841 663 665 163 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=19120 $D=1
M842 658 121 662 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=14490 $D=1
M843 659 122 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=19120 $D=1
M844 666 660 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=14490 $D=1
M845 667 661 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=19120 $D=1
M846 164 666 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=14490 $D=1
M847 657 667 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=19120 $D=1
M848 121 660 164 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=14490 $D=1
M849 122 661 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=19120 $D=1
M850 668 164 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=14490 $D=1
M851 669 657 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=19120 $D=1
M852 670 660 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=14490 $D=1
M853 671 661 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=19120 $D=1
M854 209 670 668 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=14490 $D=1
M855 210 671 669 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=19120 $D=1
M856 6 660 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=14490 $D=1
M857 7 661 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=19120 $D=1
M858 672 165 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=14490 $D=1
M859 673 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=19120 $D=1
M860 674 672 209 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=14490 $D=1
M861 675 673 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=19120 $D=1
M862 14 165 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=14490 $D=1
M863 15 165 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=19120 $D=1
M864 676 166 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=14490 $D=1
M865 677 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=19120 $D=1
M866 166 676 674 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=14490 $D=1
M867 166 677 675 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=19120 $D=1
M868 6 166 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=14490 $D=1
M869 7 166 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=19120 $D=1
M870 678 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=14490 $D=1
M871 679 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=19120 $D=1
M872 6 678 680 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=14490 $D=1
M873 7 679 681 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=19120 $D=1
M874 682 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=14490 $D=1
M875 683 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=19120 $D=1
M876 684 678 166 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=14490 $D=1
M877 685 679 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=19120 $D=1
M878 6 684 772 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=14490 $D=1
M879 7 685 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=19120 $D=1
M880 686 772 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=14490 $D=1
M881 687 773 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=19120 $D=1
M882 684 680 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=14490 $D=1
M883 685 681 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=19120 $D=1
M884 688 117 686 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=14490 $D=1
M885 689 117 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=19120 $D=1
M886 6 692 690 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=14490 $D=1
M887 7 693 691 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=19120 $D=1
M888 692 117 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=14490 $D=1
M889 693 117 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=19120 $D=1
M890 774 688 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=14490 $D=1
M891 775 689 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=19120 $D=1
M892 694 690 774 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=14490 $D=1
M893 695 691 775 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=19120 $D=1
M894 6 694 121 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=14490 $D=1
M895 7 695 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=19120 $D=1
M896 776 121 6 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=14490 $D=1
M897 777 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=19120 $D=1
M898 694 692 776 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=14490 $D=1
M899 695 693 777 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=19120 $D=1
M900 183 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=15740 $D=0
M901 184 1 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=20370 $D=0
M902 185 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=15740 $D=0
M903 186 1 3 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=20370 $D=0
M904 6 183 185 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=15740 $D=0
M905 7 184 186 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=20370 $D=0
M906 187 1 4 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=15740 $D=0
M907 188 1 4 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=20370 $D=0
M908 5 183 187 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=15740 $D=0
M909 5 184 188 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=20370 $D=0
M910 189 1 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=15740 $D=0
M911 190 1 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=20370 $D=0
M912 6 183 189 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=15740 $D=0
M913 7 184 190 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=20370 $D=0
M914 193 9 189 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=15740 $D=0
M915 194 9 190 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=20370 $D=0
M916 191 9 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=15740 $D=0
M917 192 9 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=20370 $D=0
M918 195 9 187 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=15740 $D=0
M919 196 9 188 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=20370 $D=0
M920 185 191 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=15740 $D=0
M921 186 192 196 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=20370 $D=0
M922 197 10 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=15740 $D=0
M923 198 10 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=20370 $D=0
M924 199 10 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=15740 $D=0
M925 200 10 196 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=20370 $D=0
M926 193 197 199 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=15740 $D=0
M927 194 198 200 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=20370 $D=0
M928 201 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=15740 $D=0
M929 202 11 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=20370 $D=0
M930 203 11 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=15740 $D=0
M931 204 11 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=20370 $D=0
M932 12 201 203 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=15740 $D=0
M933 13 202 204 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=20370 $D=0
M934 205 11 14 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=15740 $D=0
M935 206 11 15 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=20370 $D=0
M936 207 201 205 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=15740 $D=0
M937 208 202 206 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=20370 $D=0
M938 211 11 209 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=15740 $D=0
M939 212 11 210 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=20370 $D=0
M940 199 201 211 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=15740 $D=0
M941 200 202 212 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=20370 $D=0
M942 215 16 211 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=15740 $D=0
M943 216 16 212 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=20370 $D=0
M944 213 16 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=15740 $D=0
M945 214 16 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=20370 $D=0
M946 217 16 205 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=15740 $D=0
M947 218 16 206 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=20370 $D=0
M948 203 213 217 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=15740 $D=0
M949 204 214 218 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=20370 $D=0
M950 219 17 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=15740 $D=0
M951 220 17 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=20370 $D=0
M952 221 17 217 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=15740 $D=0
M953 222 17 218 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=20370 $D=0
M954 215 219 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=15740 $D=0
M955 216 220 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=20370 $D=0
M956 167 18 223 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=15740 $D=0
M957 168 18 224 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=20370 $D=0
M958 225 19 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=15740 $D=0
M959 226 19 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=20370 $D=0
M960 227 223 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=15740 $D=0
M961 228 224 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=20370 $D=0
M962 167 227 696 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=15740 $D=0
M963 168 228 697 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=20370 $D=0
M964 229 696 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=15740 $D=0
M965 230 697 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=20370 $D=0
M966 227 18 229 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=15740 $D=0
M967 228 18 230 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=20370 $D=0
M968 229 225 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=15740 $D=0
M969 230 226 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=20370 $D=0
M970 235 233 229 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=15740 $D=0
M971 236 234 230 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=20370 $D=0
M972 233 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=15740 $D=0
M973 234 20 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=20370 $D=0
M974 167 21 237 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=15740 $D=0
M975 168 21 238 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=20370 $D=0
M976 239 22 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=15740 $D=0
M977 240 22 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=20370 $D=0
M978 241 237 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=15740 $D=0
M979 242 238 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=20370 $D=0
M980 167 241 698 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=15740 $D=0
M981 168 242 699 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=20370 $D=0
M982 243 698 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=15740 $D=0
M983 244 699 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=20370 $D=0
M984 241 21 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=15740 $D=0
M985 242 21 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=20370 $D=0
M986 243 239 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=15740 $D=0
M987 244 240 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=20370 $D=0
M988 235 245 243 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=15740 $D=0
M989 236 246 244 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=20370 $D=0
M990 245 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=15740 $D=0
M991 246 23 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=20370 $D=0
M992 167 24 247 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=15740 $D=0
M993 168 24 248 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=20370 $D=0
M994 249 25 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=15740 $D=0
M995 250 25 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=20370 $D=0
M996 251 247 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=15740 $D=0
M997 252 248 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=20370 $D=0
M998 167 251 700 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=15740 $D=0
M999 168 252 701 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=20370 $D=0
M1000 253 700 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=15740 $D=0
M1001 254 701 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=20370 $D=0
M1002 251 24 253 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=15740 $D=0
M1003 252 24 254 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=20370 $D=0
M1004 253 249 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=15740 $D=0
M1005 254 250 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=20370 $D=0
M1006 235 255 253 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=15740 $D=0
M1007 236 256 254 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=20370 $D=0
M1008 255 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=15740 $D=0
M1009 256 26 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=20370 $D=0
M1010 167 27 257 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=15740 $D=0
M1011 168 27 258 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=20370 $D=0
M1012 259 28 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=15740 $D=0
M1013 260 28 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=20370 $D=0
M1014 261 257 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=15740 $D=0
M1015 262 258 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=20370 $D=0
M1016 167 261 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=15740 $D=0
M1017 168 262 703 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=20370 $D=0
M1018 263 702 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=15740 $D=0
M1019 264 703 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=20370 $D=0
M1020 261 27 263 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=15740 $D=0
M1021 262 27 264 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=20370 $D=0
M1022 263 259 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=15740 $D=0
M1023 264 260 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=20370 $D=0
M1024 235 265 263 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=15740 $D=0
M1025 236 266 264 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=20370 $D=0
M1026 265 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=15740 $D=0
M1027 266 29 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=20370 $D=0
M1028 167 30 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=15740 $D=0
M1029 168 30 268 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=20370 $D=0
M1030 269 31 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=15740 $D=0
M1031 270 31 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=20370 $D=0
M1032 271 267 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=15740 $D=0
M1033 272 268 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=20370 $D=0
M1034 167 271 704 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=15740 $D=0
M1035 168 272 705 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=20370 $D=0
M1036 273 704 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=15740 $D=0
M1037 274 705 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=20370 $D=0
M1038 271 30 273 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=15740 $D=0
M1039 272 30 274 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=20370 $D=0
M1040 273 269 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=15740 $D=0
M1041 274 270 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=20370 $D=0
M1042 235 275 273 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=15740 $D=0
M1043 236 276 274 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=20370 $D=0
M1044 275 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=15740 $D=0
M1045 276 32 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=20370 $D=0
M1046 167 33 277 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=15740 $D=0
M1047 168 33 278 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=20370 $D=0
M1048 279 34 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=15740 $D=0
M1049 280 34 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=20370 $D=0
M1050 281 277 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=15740 $D=0
M1051 282 278 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=20370 $D=0
M1052 167 281 706 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=15740 $D=0
M1053 168 282 707 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=20370 $D=0
M1054 283 706 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=15740 $D=0
M1055 284 707 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=20370 $D=0
M1056 281 33 283 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=15740 $D=0
M1057 282 33 284 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=20370 $D=0
M1058 283 279 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=15740 $D=0
M1059 284 280 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=20370 $D=0
M1060 235 285 283 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=15740 $D=0
M1061 236 286 284 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=20370 $D=0
M1062 285 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=15740 $D=0
M1063 286 35 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=20370 $D=0
M1064 167 36 287 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=15740 $D=0
M1065 168 36 288 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=20370 $D=0
M1066 289 37 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=15740 $D=0
M1067 290 37 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=20370 $D=0
M1068 291 287 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=15740 $D=0
M1069 292 288 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=20370 $D=0
M1070 167 291 708 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=15740 $D=0
M1071 168 292 709 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=20370 $D=0
M1072 293 708 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=15740 $D=0
M1073 294 709 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=20370 $D=0
M1074 291 36 293 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=15740 $D=0
M1075 292 36 294 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=20370 $D=0
M1076 293 289 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=15740 $D=0
M1077 294 290 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=20370 $D=0
M1078 235 295 293 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=15740 $D=0
M1079 236 296 294 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=20370 $D=0
M1080 295 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=15740 $D=0
M1081 296 38 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=20370 $D=0
M1082 167 39 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=15740 $D=0
M1083 168 39 298 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=20370 $D=0
M1084 299 40 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=15740 $D=0
M1085 300 40 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=20370 $D=0
M1086 301 297 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=15740 $D=0
M1087 302 298 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=20370 $D=0
M1088 167 301 710 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=15740 $D=0
M1089 168 302 711 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=20370 $D=0
M1090 303 710 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=15740 $D=0
M1091 304 711 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=20370 $D=0
M1092 301 39 303 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=15740 $D=0
M1093 302 39 304 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=20370 $D=0
M1094 303 299 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=15740 $D=0
M1095 304 300 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=20370 $D=0
M1096 235 305 303 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=15740 $D=0
M1097 236 306 304 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=20370 $D=0
M1098 305 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=15740 $D=0
M1099 306 41 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=20370 $D=0
M1100 167 42 307 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=15740 $D=0
M1101 168 42 308 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=20370 $D=0
M1102 309 43 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=15740 $D=0
M1103 310 43 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=20370 $D=0
M1104 311 307 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=15740 $D=0
M1105 312 308 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=20370 $D=0
M1106 167 311 712 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=15740 $D=0
M1107 168 312 713 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=20370 $D=0
M1108 313 712 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=15740 $D=0
M1109 314 713 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=20370 $D=0
M1110 311 42 313 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=15740 $D=0
M1111 312 42 314 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=20370 $D=0
M1112 313 309 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=15740 $D=0
M1113 314 310 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=20370 $D=0
M1114 235 315 313 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=15740 $D=0
M1115 236 316 314 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=20370 $D=0
M1116 315 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=15740 $D=0
M1117 316 44 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=20370 $D=0
M1118 167 45 317 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=15740 $D=0
M1119 168 45 318 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=20370 $D=0
M1120 319 46 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=15740 $D=0
M1121 320 46 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=20370 $D=0
M1122 321 317 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=15740 $D=0
M1123 322 318 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=20370 $D=0
M1124 167 321 714 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=15740 $D=0
M1125 168 322 715 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=20370 $D=0
M1126 323 714 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=15740 $D=0
M1127 324 715 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=20370 $D=0
M1128 321 45 323 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=15740 $D=0
M1129 322 45 324 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=20370 $D=0
M1130 323 319 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=15740 $D=0
M1131 324 320 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=20370 $D=0
M1132 235 325 323 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=15740 $D=0
M1133 236 326 324 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=20370 $D=0
M1134 325 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=15740 $D=0
M1135 326 47 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=20370 $D=0
M1136 167 48 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=15740 $D=0
M1137 168 48 328 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=20370 $D=0
M1138 329 49 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=15740 $D=0
M1139 330 49 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=20370 $D=0
M1140 331 327 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=15740 $D=0
M1141 332 328 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=20370 $D=0
M1142 167 331 716 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=15740 $D=0
M1143 168 332 717 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=20370 $D=0
M1144 333 716 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=15740 $D=0
M1145 334 717 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=20370 $D=0
M1146 331 48 333 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=15740 $D=0
M1147 332 48 334 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=20370 $D=0
M1148 333 329 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=15740 $D=0
M1149 334 330 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=20370 $D=0
M1150 235 335 333 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=15740 $D=0
M1151 236 336 334 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=20370 $D=0
M1152 335 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=15740 $D=0
M1153 336 50 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=20370 $D=0
M1154 167 51 337 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=15740 $D=0
M1155 168 51 338 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=20370 $D=0
M1156 339 52 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=15740 $D=0
M1157 340 52 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=20370 $D=0
M1158 341 337 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=15740 $D=0
M1159 342 338 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=20370 $D=0
M1160 167 341 718 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=15740 $D=0
M1161 168 342 719 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=20370 $D=0
M1162 343 718 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=15740 $D=0
M1163 344 719 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=20370 $D=0
M1164 341 51 343 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=15740 $D=0
M1165 342 51 344 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=20370 $D=0
M1166 343 339 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=15740 $D=0
M1167 344 340 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=20370 $D=0
M1168 235 345 343 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=15740 $D=0
M1169 236 346 344 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=20370 $D=0
M1170 345 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=15740 $D=0
M1171 346 53 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=20370 $D=0
M1172 167 54 347 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=15740 $D=0
M1173 168 54 348 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=20370 $D=0
M1174 349 55 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=15740 $D=0
M1175 350 55 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=20370 $D=0
M1176 351 347 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=15740 $D=0
M1177 352 348 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=20370 $D=0
M1178 167 351 720 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=15740 $D=0
M1179 168 352 721 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=20370 $D=0
M1180 353 720 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=15740 $D=0
M1181 354 721 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=20370 $D=0
M1182 351 54 353 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=15740 $D=0
M1183 352 54 354 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=20370 $D=0
M1184 353 349 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=15740 $D=0
M1185 354 350 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=20370 $D=0
M1186 235 355 353 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=15740 $D=0
M1187 236 356 354 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=20370 $D=0
M1188 355 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=15740 $D=0
M1189 356 56 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=20370 $D=0
M1190 167 57 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=15740 $D=0
M1191 168 57 358 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=20370 $D=0
M1192 359 58 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=15740 $D=0
M1193 360 58 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=20370 $D=0
M1194 361 357 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=15740 $D=0
M1195 362 358 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=20370 $D=0
M1196 167 361 722 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=15740 $D=0
M1197 168 362 723 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=20370 $D=0
M1198 363 722 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=15740 $D=0
M1199 364 723 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=20370 $D=0
M1200 361 57 363 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=15740 $D=0
M1201 362 57 364 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=20370 $D=0
M1202 363 359 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=15740 $D=0
M1203 364 360 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=20370 $D=0
M1204 235 365 363 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=15740 $D=0
M1205 236 366 364 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=20370 $D=0
M1206 365 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=15740 $D=0
M1207 366 59 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=20370 $D=0
M1208 167 60 367 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=15740 $D=0
M1209 168 60 368 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=20370 $D=0
M1210 369 61 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=15740 $D=0
M1211 370 61 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=20370 $D=0
M1212 371 367 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=15740 $D=0
M1213 372 368 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=20370 $D=0
M1214 167 371 724 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=15740 $D=0
M1215 168 372 725 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=20370 $D=0
M1216 373 724 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=15740 $D=0
M1217 374 725 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=20370 $D=0
M1218 371 60 373 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=15740 $D=0
M1219 372 60 374 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=20370 $D=0
M1220 373 369 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=15740 $D=0
M1221 374 370 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=20370 $D=0
M1222 235 375 373 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=15740 $D=0
M1223 236 376 374 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=20370 $D=0
M1224 375 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=15740 $D=0
M1225 376 62 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=20370 $D=0
M1226 167 63 377 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=15740 $D=0
M1227 168 63 378 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=20370 $D=0
M1228 379 64 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=15740 $D=0
M1229 380 64 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=20370 $D=0
M1230 381 377 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=15740 $D=0
M1231 382 378 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=20370 $D=0
M1232 167 381 726 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=15740 $D=0
M1233 168 382 727 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=20370 $D=0
M1234 383 726 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=15740 $D=0
M1235 384 727 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=20370 $D=0
M1236 381 63 383 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=15740 $D=0
M1237 382 63 384 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=20370 $D=0
M1238 383 379 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=15740 $D=0
M1239 384 380 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=20370 $D=0
M1240 235 385 383 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=15740 $D=0
M1241 236 386 384 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=20370 $D=0
M1242 385 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=15740 $D=0
M1243 386 65 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=20370 $D=0
M1244 167 66 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=15740 $D=0
M1245 168 66 388 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=20370 $D=0
M1246 389 67 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=15740 $D=0
M1247 390 67 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=20370 $D=0
M1248 391 387 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=15740 $D=0
M1249 392 388 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=20370 $D=0
M1250 167 391 728 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=15740 $D=0
M1251 168 392 729 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=20370 $D=0
M1252 393 728 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=15740 $D=0
M1253 394 729 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=20370 $D=0
M1254 391 66 393 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=15740 $D=0
M1255 392 66 394 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=20370 $D=0
M1256 393 389 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=15740 $D=0
M1257 394 390 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=20370 $D=0
M1258 235 395 393 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=15740 $D=0
M1259 236 396 394 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=20370 $D=0
M1260 395 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=15740 $D=0
M1261 396 68 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=20370 $D=0
M1262 167 69 397 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=15740 $D=0
M1263 168 69 398 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=20370 $D=0
M1264 399 70 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=15740 $D=0
M1265 400 70 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=20370 $D=0
M1266 401 397 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=15740 $D=0
M1267 402 398 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=20370 $D=0
M1268 167 401 730 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=15740 $D=0
M1269 168 402 731 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=20370 $D=0
M1270 403 730 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=15740 $D=0
M1271 404 731 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=20370 $D=0
M1272 401 69 403 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=15740 $D=0
M1273 402 69 404 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=20370 $D=0
M1274 403 399 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=15740 $D=0
M1275 404 400 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=20370 $D=0
M1276 235 405 403 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=15740 $D=0
M1277 236 406 404 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=20370 $D=0
M1278 405 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=15740 $D=0
M1279 406 71 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=20370 $D=0
M1280 167 72 407 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=15740 $D=0
M1281 168 72 408 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=20370 $D=0
M1282 409 73 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=15740 $D=0
M1283 410 73 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=20370 $D=0
M1284 411 407 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=15740 $D=0
M1285 412 408 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=20370 $D=0
M1286 167 411 732 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=15740 $D=0
M1287 168 412 733 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=20370 $D=0
M1288 413 732 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=15740 $D=0
M1289 414 733 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=20370 $D=0
M1290 411 72 413 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=15740 $D=0
M1291 412 72 414 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=20370 $D=0
M1292 413 409 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=15740 $D=0
M1293 414 410 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=20370 $D=0
M1294 235 415 413 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=15740 $D=0
M1295 236 416 414 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=20370 $D=0
M1296 415 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=15740 $D=0
M1297 416 74 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=20370 $D=0
M1298 167 75 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=15740 $D=0
M1299 168 75 418 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=20370 $D=0
M1300 419 76 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=15740 $D=0
M1301 420 76 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=20370 $D=0
M1302 421 417 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=15740 $D=0
M1303 422 418 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=20370 $D=0
M1304 167 421 734 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=15740 $D=0
M1305 168 422 735 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=20370 $D=0
M1306 423 734 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=15740 $D=0
M1307 424 735 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=20370 $D=0
M1308 421 75 423 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=15740 $D=0
M1309 422 75 424 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=20370 $D=0
M1310 423 419 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=15740 $D=0
M1311 424 420 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=20370 $D=0
M1312 235 425 423 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=15740 $D=0
M1313 236 426 424 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=20370 $D=0
M1314 425 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=15740 $D=0
M1315 426 77 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=20370 $D=0
M1316 167 78 427 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=15740 $D=0
M1317 168 78 428 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=20370 $D=0
M1318 429 79 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=15740 $D=0
M1319 430 79 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=20370 $D=0
M1320 431 427 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=15740 $D=0
M1321 432 428 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=20370 $D=0
M1322 167 431 736 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=15740 $D=0
M1323 168 432 737 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=20370 $D=0
M1324 433 736 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=15740 $D=0
M1325 434 737 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=20370 $D=0
M1326 431 78 433 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=15740 $D=0
M1327 432 78 434 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=20370 $D=0
M1328 433 429 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=15740 $D=0
M1329 434 430 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=20370 $D=0
M1330 235 435 433 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=15740 $D=0
M1331 236 436 434 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=20370 $D=0
M1332 435 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=15740 $D=0
M1333 436 80 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=20370 $D=0
M1334 167 81 437 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=15740 $D=0
M1335 168 81 438 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=20370 $D=0
M1336 439 82 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=15740 $D=0
M1337 440 82 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=20370 $D=0
M1338 441 437 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=15740 $D=0
M1339 442 438 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=20370 $D=0
M1340 167 441 738 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=15740 $D=0
M1341 168 442 739 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=20370 $D=0
M1342 443 738 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=15740 $D=0
M1343 444 739 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=20370 $D=0
M1344 441 81 443 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=15740 $D=0
M1345 442 81 444 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=20370 $D=0
M1346 443 439 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=15740 $D=0
M1347 444 440 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=20370 $D=0
M1348 235 445 443 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=15740 $D=0
M1349 236 446 444 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=20370 $D=0
M1350 445 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=15740 $D=0
M1351 446 83 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=20370 $D=0
M1352 167 84 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=15740 $D=0
M1353 168 84 448 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=20370 $D=0
M1354 449 85 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=15740 $D=0
M1355 450 85 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=20370 $D=0
M1356 451 447 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=15740 $D=0
M1357 452 448 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=20370 $D=0
M1358 167 451 740 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=15740 $D=0
M1359 168 452 741 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=20370 $D=0
M1360 453 740 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=15740 $D=0
M1361 454 741 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=20370 $D=0
M1362 451 84 453 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=15740 $D=0
M1363 452 84 454 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=20370 $D=0
M1364 453 449 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=15740 $D=0
M1365 454 450 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=20370 $D=0
M1366 235 455 453 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=15740 $D=0
M1367 236 456 454 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=20370 $D=0
M1368 455 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=15740 $D=0
M1369 456 86 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=20370 $D=0
M1370 167 87 457 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=15740 $D=0
M1371 168 87 458 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=20370 $D=0
M1372 459 88 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=15740 $D=0
M1373 460 88 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=20370 $D=0
M1374 461 457 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=15740 $D=0
M1375 462 458 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=20370 $D=0
M1376 167 461 742 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=15740 $D=0
M1377 168 462 743 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=20370 $D=0
M1378 463 742 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=15740 $D=0
M1379 464 743 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=20370 $D=0
M1380 461 87 463 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=15740 $D=0
M1381 462 87 464 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=20370 $D=0
M1382 463 459 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=15740 $D=0
M1383 464 460 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=20370 $D=0
M1384 235 465 463 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=15740 $D=0
M1385 236 466 464 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=20370 $D=0
M1386 465 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=15740 $D=0
M1387 466 89 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=20370 $D=0
M1388 167 90 467 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=15740 $D=0
M1389 168 90 468 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=20370 $D=0
M1390 469 91 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=15740 $D=0
M1391 470 91 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=20370 $D=0
M1392 471 467 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=15740 $D=0
M1393 472 468 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=20370 $D=0
M1394 167 471 744 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=15740 $D=0
M1395 168 472 745 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=20370 $D=0
M1396 473 744 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=15740 $D=0
M1397 474 745 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=20370 $D=0
M1398 471 90 473 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=15740 $D=0
M1399 472 90 474 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=20370 $D=0
M1400 473 469 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=15740 $D=0
M1401 474 470 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=20370 $D=0
M1402 235 475 473 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=15740 $D=0
M1403 236 476 474 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=20370 $D=0
M1404 475 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=15740 $D=0
M1405 476 92 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=20370 $D=0
M1406 167 93 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=15740 $D=0
M1407 168 93 478 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=20370 $D=0
M1408 479 94 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=15740 $D=0
M1409 480 94 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=20370 $D=0
M1410 481 477 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=15740 $D=0
M1411 482 478 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=20370 $D=0
M1412 167 481 746 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=15740 $D=0
M1413 168 482 747 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=20370 $D=0
M1414 483 746 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=15740 $D=0
M1415 484 747 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=20370 $D=0
M1416 481 93 483 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=15740 $D=0
M1417 482 93 484 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=20370 $D=0
M1418 483 479 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=15740 $D=0
M1419 484 480 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=20370 $D=0
M1420 235 485 483 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=15740 $D=0
M1421 236 486 484 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=20370 $D=0
M1422 485 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=15740 $D=0
M1423 486 95 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=20370 $D=0
M1424 167 96 487 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=15740 $D=0
M1425 168 96 488 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=20370 $D=0
M1426 489 97 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=15740 $D=0
M1427 490 97 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=20370 $D=0
M1428 491 487 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=15740 $D=0
M1429 492 488 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=20370 $D=0
M1430 167 491 748 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=15740 $D=0
M1431 168 492 749 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=20370 $D=0
M1432 493 748 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=15740 $D=0
M1433 494 749 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=20370 $D=0
M1434 491 96 493 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=15740 $D=0
M1435 492 96 494 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=20370 $D=0
M1436 493 489 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=15740 $D=0
M1437 494 490 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=20370 $D=0
M1438 235 495 493 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=15740 $D=0
M1439 236 496 494 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=20370 $D=0
M1440 495 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=15740 $D=0
M1441 496 98 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=20370 $D=0
M1442 167 99 497 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=15740 $D=0
M1443 168 99 498 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=20370 $D=0
M1444 499 100 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=15740 $D=0
M1445 500 100 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=20370 $D=0
M1446 501 497 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=15740 $D=0
M1447 502 498 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=20370 $D=0
M1448 167 501 750 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=15740 $D=0
M1449 168 502 751 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=20370 $D=0
M1450 503 750 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=15740 $D=0
M1451 504 751 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=20370 $D=0
M1452 501 99 503 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=15740 $D=0
M1453 502 99 504 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=20370 $D=0
M1454 503 499 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=15740 $D=0
M1455 504 500 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=20370 $D=0
M1456 235 505 503 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=15740 $D=0
M1457 236 506 504 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=20370 $D=0
M1458 505 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=15740 $D=0
M1459 506 101 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=20370 $D=0
M1460 167 102 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=15740 $D=0
M1461 168 102 508 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=20370 $D=0
M1462 509 103 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=15740 $D=0
M1463 510 103 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=20370 $D=0
M1464 511 507 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=15740 $D=0
M1465 512 508 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=20370 $D=0
M1466 167 511 752 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=15740 $D=0
M1467 168 512 753 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=20370 $D=0
M1468 513 752 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=15740 $D=0
M1469 514 753 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=20370 $D=0
M1470 511 102 513 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=15740 $D=0
M1471 512 102 514 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=20370 $D=0
M1472 513 509 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=15740 $D=0
M1473 514 510 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=20370 $D=0
M1474 235 515 513 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=15740 $D=0
M1475 236 516 514 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=20370 $D=0
M1476 515 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=15740 $D=0
M1477 516 104 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=20370 $D=0
M1478 167 105 517 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=15740 $D=0
M1479 168 105 518 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=20370 $D=0
M1480 519 106 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=15740 $D=0
M1481 520 106 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=20370 $D=0
M1482 521 517 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=15740 $D=0
M1483 522 518 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=20370 $D=0
M1484 167 521 754 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=15740 $D=0
M1485 168 522 755 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=20370 $D=0
M1486 523 754 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=15740 $D=0
M1487 524 755 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=20370 $D=0
M1488 521 105 523 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=15740 $D=0
M1489 522 105 524 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=20370 $D=0
M1490 523 519 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=15740 $D=0
M1491 524 520 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=20370 $D=0
M1492 235 525 523 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=15740 $D=0
M1493 236 526 524 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=20370 $D=0
M1494 525 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=15740 $D=0
M1495 526 108 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=20370 $D=0
M1496 167 110 527 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=15740 $D=0
M1497 168 110 528 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=20370 $D=0
M1498 529 111 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=15740 $D=0
M1499 530 111 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=20370 $D=0
M1500 531 527 221 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=15740 $D=0
M1501 532 528 222 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=20370 $D=0
M1502 167 531 756 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=15740 $D=0
M1503 168 532 757 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=20370 $D=0
M1504 533 756 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=15740 $D=0
M1505 534 757 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=20370 $D=0
M1506 531 110 533 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=15740 $D=0
M1507 532 110 534 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=20370 $D=0
M1508 533 529 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=15740 $D=0
M1509 534 530 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=20370 $D=0
M1510 235 535 533 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=15740 $D=0
M1511 236 536 534 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=20370 $D=0
M1512 535 114 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=15740 $D=0
M1513 536 114 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=20370 $D=0
M1514 167 115 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=15740 $D=0
M1515 168 115 538 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=20370 $D=0
M1516 539 116 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=15740 $D=0
M1517 540 116 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=20370 $D=0
M1518 6 539 231 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=15740 $D=0
M1519 7 540 232 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=20370 $D=0
M1520 235 537 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=15740 $D=0
M1521 236 538 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=20370 $D=0
M1522 167 543 541 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=15740 $D=0
M1523 168 544 542 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=20370 $D=0
M1524 543 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=15740 $D=0
M1525 544 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=20370 $D=0
M1526 758 231 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=15740 $D=0
M1527 759 232 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=20370 $D=0
M1528 545 543 758 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=15740 $D=0
M1529 546 544 759 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=20370 $D=0
M1530 167 545 547 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=15740 $D=0
M1531 168 546 548 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=20370 $D=0
M1532 760 547 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=15740 $D=0
M1533 761 548 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=20370 $D=0
M1534 545 541 760 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=15740 $D=0
M1535 546 542 761 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=20370 $D=0
M1536 167 551 549 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=15740 $D=0
M1537 168 552 550 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=20370 $D=0
M1538 551 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=15740 $D=0
M1539 552 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=20370 $D=0
M1540 762 235 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=15740 $D=0
M1541 763 236 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=20370 $D=0
M1542 553 551 762 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=15740 $D=0
M1543 554 552 763 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=20370 $D=0
M1544 167 553 118 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=15740 $D=0
M1545 168 554 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=20370 $D=0
M1546 764 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=15740 $D=0
M1547 765 119 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=20370 $D=0
M1548 553 549 764 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=15740 $D=0
M1549 554 550 765 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=20370 $D=0
M1550 555 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=15740 $D=0
M1551 556 120 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=20370 $D=0
M1552 557 120 547 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=15740 $D=0
M1553 558 120 548 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=20370 $D=0
M1554 121 555 557 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=15740 $D=0
M1555 122 556 558 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=20370 $D=0
M1556 559 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=15740 $D=0
M1557 560 123 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=20370 $D=0
M1558 562 123 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=15740 $D=0
M1559 563 123 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=20370 $D=0
M1560 766 559 562 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=15740 $D=0
M1561 767 560 563 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=20370 $D=0
M1562 167 561 766 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=15740 $D=0
M1563 168 119 767 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=20370 $D=0
M1564 564 124 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=15740 $D=0
M1565 565 124 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=20370 $D=0
M1566 566 124 562 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=15740 $D=0
M1567 567 124 563 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=20370 $D=0
M1568 12 564 566 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=15740 $D=0
M1569 13 565 567 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=20370 $D=0
M1570 569 568 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=15740 $D=0
M1571 570 125 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=20370 $D=0
M1572 167 573 571 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=15740 $D=0
M1573 168 574 572 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=20370 $D=0
M1574 575 557 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=15740 $D=0
M1575 576 558 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=20370 $D=0
M1576 573 557 568 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=15740 $D=0
M1577 574 558 125 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=20370 $D=0
M1578 569 575 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=15740 $D=0
M1579 570 576 574 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=20370 $D=0
M1580 577 571 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=15740 $D=0
M1581 578 572 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=20370 $D=0
M1582 126 571 566 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=15740 $D=0
M1583 568 572 567 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=20370 $D=0
M1584 557 577 126 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=15740 $D=0
M1585 558 578 568 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=20370 $D=0
M1586 579 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=15740 $D=0
M1587 580 568 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=20370 $D=0
M1588 581 571 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=15740 $D=0
M1589 582 572 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=20370 $D=0
M1590 583 571 579 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=15740 $D=0
M1591 584 572 580 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=20370 $D=0
M1592 566 581 583 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=15740 $D=0
M1593 567 582 584 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=20370 $D=0
M1594 778 557 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=15380 $D=0
M1595 779 558 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=20010 $D=0
M1596 585 566 778 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=15380 $D=0
M1597 586 567 779 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=20010 $D=0
M1598 587 583 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=15740 $D=0
M1599 588 584 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=20370 $D=0
M1600 589 557 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=15740 $D=0
M1601 590 558 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=20370 $D=0
M1602 167 566 589 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=15740 $D=0
M1603 168 567 590 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=20370 $D=0
M1604 591 557 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=15740 $D=0
M1605 592 558 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=20370 $D=0
M1606 167 566 591 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=15740 $D=0
M1607 168 567 592 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=20370 $D=0
M1608 780 557 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=15560 $D=0
M1609 781 558 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=20190 $D=0
M1610 595 566 780 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=15560 $D=0
M1611 596 567 781 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=20190 $D=0
M1612 167 591 595 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=15740 $D=0
M1613 168 592 596 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=20370 $D=0
M1614 597 129 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=15740 $D=0
M1615 598 129 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=20370 $D=0
M1616 599 129 585 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=15740 $D=0
M1617 600 129 586 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=20370 $D=0
M1618 589 597 599 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=15740 $D=0
M1619 590 598 600 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=20370 $D=0
M1620 601 129 587 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=15740 $D=0
M1621 602 129 588 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=20370 $D=0
M1622 595 597 601 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=15740 $D=0
M1623 596 598 602 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=20370 $D=0
M1624 603 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=15740 $D=0
M1625 604 130 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=20370 $D=0
M1626 605 130 601 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=15740 $D=0
M1627 606 130 602 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=20370 $D=0
M1628 599 603 605 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=15740 $D=0
M1629 600 604 606 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=20370 $D=0
M1630 14 605 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=15740 $D=0
M1631 15 606 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=20370 $D=0
M1632 607 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=15740 $D=0
M1633 608 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=20370 $D=0
M1634 609 131 132 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=15740 $D=0
M1635 610 131 133 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=20370 $D=0
M1636 134 607 609 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=15740 $D=0
M1637 135 608 610 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=20370 $D=0
M1638 611 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=15740 $D=0
M1639 612 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=20370 $D=0
M1640 613 131 136 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=15740 $D=0
M1641 614 131 137 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=20370 $D=0
M1642 138 611 613 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=15740 $D=0
M1643 139 612 614 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=20370 $D=0
M1644 615 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=15740 $D=0
M1645 616 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=20370 $D=0
M1646 617 131 127 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=15740 $D=0
M1647 618 131 128 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=20370 $D=0
M1648 140 615 617 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=15740 $D=0
M1649 141 616 618 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=20370 $D=0
M1650 619 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=15740 $D=0
M1651 620 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=20370 $D=0
M1652 621 131 143 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=15740 $D=0
M1653 622 131 144 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=20370 $D=0
M1654 140 619 621 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=15740 $D=0
M1655 140 620 622 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=20370 $D=0
M1656 623 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=15740 $D=0
M1657 624 131 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=20370 $D=0
M1658 625 131 145 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=15740 $D=0
M1659 626 131 146 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=20370 $D=0
M1660 140 623 625 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=15740 $D=0
M1661 140 624 626 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=20370 $D=0
M1662 167 557 768 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=15740 $D=0
M1663 168 558 769 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=20370 $D=0
M1664 135 768 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=15740 $D=0
M1665 132 769 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=20370 $D=0
M1666 627 147 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=15740 $D=0
M1667 628 147 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=20370 $D=0
M1668 148 147 135 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=15740 $D=0
M1669 149 147 132 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=20370 $D=0
M1670 609 627 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=15740 $D=0
M1671 610 628 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=20370 $D=0
M1672 629 150 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=15740 $D=0
M1673 630 150 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=20370 $D=0
M1674 151 150 148 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=15740 $D=0
M1675 107 150 149 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=20370 $D=0
M1676 613 629 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=15740 $D=0
M1677 614 630 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=20370 $D=0
M1678 631 152 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=15740 $D=0
M1679 632 152 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=20370 $D=0
M1680 153 152 151 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=15740 $D=0
M1681 112 152 107 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=20370 $D=0
M1682 617 631 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=15740 $D=0
M1683 618 632 112 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=20370 $D=0
M1684 633 154 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=15740 $D=0
M1685 634 154 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=20370 $D=0
M1686 155 154 153 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=15740 $D=0
M1687 156 154 112 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=20370 $D=0
M1688 621 633 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=15740 $D=0
M1689 622 634 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=20370 $D=0
M1690 635 157 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=15740 $D=0
M1691 636 157 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=20370 $D=0
M1692 207 157 155 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=15740 $D=0
M1693 208 157 156 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=20370 $D=0
M1694 625 635 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=15740 $D=0
M1695 626 636 208 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=20370 $D=0
M1696 637 158 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=15740 $D=0
M1697 638 158 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=20370 $D=0
M1698 639 158 561 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=15740 $D=0
M1699 640 158 119 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=20370 $D=0
M1700 12 637 639 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=15740 $D=0
M1701 13 638 640 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=20370 $D=0
M1702 641 547 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=15740 $D=0
M1703 642 548 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=20370 $D=0
M1704 167 639 641 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=15740 $D=0
M1705 168 640 642 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=20370 $D=0
M1706 782 547 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=15560 $D=0
M1707 783 548 168 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=20190 $D=0
M1708 645 639 782 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=15560 $D=0
M1709 646 640 783 168 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=20190 $D=0
M1710 167 641 645 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=15740 $D=0
M1711 168 642 646 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=20370 $D=0
M1712 770 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=15740 $D=0
M1713 771 647 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=20370 $D=0
M1714 167 645 770 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=15740 $D=0
M1715 168 646 771 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=20370 $D=0
M1716 647 770 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=15740 $D=0
M1717 160 771 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=20370 $D=0
M1718 784 547 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=15380 $D=0
M1719 785 548 168 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=20010 $D=0
M1720 648 650 784 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=15380 $D=0
M1721 649 651 785 168 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=20010 $D=0
M1722 650 639 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=15740 $D=0
M1723 651 640 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=20370 $D=0
M1724 652 648 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=15740 $D=0
M1725 653 649 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=20370 $D=0
M1726 167 159 652 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=15740 $D=0
M1727 168 647 653 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=20370 $D=0
M1728 655 161 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=15740 $D=0
M1729 656 654 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=20370 $D=0
M1730 654 652 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=15740 $D=0
M1731 162 653 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=20370 $D=0
M1732 167 655 654 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=15740 $D=0
M1733 168 656 162 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=20370 $D=0
M1734 658 657 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=15740 $D=0
M1735 659 163 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=20370 $D=0
M1736 167 662 660 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=15740 $D=0
M1737 168 663 661 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=20370 $D=0
M1738 664 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=15740 $D=0
M1739 665 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=20370 $D=0
M1740 662 121 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=15740 $D=0
M1741 663 122 163 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=20370 $D=0
M1742 658 664 662 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=15740 $D=0
M1743 659 665 663 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=20370 $D=0
M1744 666 660 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=15740 $D=0
M1745 667 661 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=20370 $D=0
M1746 164 660 6 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=15740 $D=0
M1747 657 661 7 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=20370 $D=0
M1748 121 666 164 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=15740 $D=0
M1749 122 667 657 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=20370 $D=0
M1750 668 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=15740 $D=0
M1751 669 657 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=20370 $D=0
M1752 670 660 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=15740 $D=0
M1753 671 661 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=20370 $D=0
M1754 209 660 668 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=15740 $D=0
M1755 210 661 669 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=20370 $D=0
M1756 6 670 209 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=15740 $D=0
M1757 7 671 210 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=20370 $D=0
M1758 672 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=15740 $D=0
M1759 673 165 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=20370 $D=0
M1760 674 165 209 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=15740 $D=0
M1761 675 165 210 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=20370 $D=0
M1762 14 672 674 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=15740 $D=0
M1763 15 673 675 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=20370 $D=0
M1764 676 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=15740 $D=0
M1765 677 166 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=20370 $D=0
M1766 166 166 674 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=15740 $D=0
M1767 166 166 675 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=20370 $D=0
M1768 6 676 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=15740 $D=0
M1769 7 677 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=20370 $D=0
M1770 678 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=15740 $D=0
M1771 679 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=20370 $D=0
M1772 167 678 680 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=15740 $D=0
M1773 168 679 681 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=20370 $D=0
M1774 682 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=15740 $D=0
M1775 683 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=20370 $D=0
M1776 684 680 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=15740 $D=0
M1777 685 681 166 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=20370 $D=0
M1778 167 684 772 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=15740 $D=0
M1779 168 685 773 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=20370 $D=0
M1780 686 772 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=15740 $D=0
M1781 687 773 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=20370 $D=0
M1782 684 678 686 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=15740 $D=0
M1783 685 679 687 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=20370 $D=0
M1784 688 682 686 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=15740 $D=0
M1785 689 683 687 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=20370 $D=0
M1786 167 692 690 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=15740 $D=0
M1787 168 693 691 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=20370 $D=0
M1788 692 117 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=15740 $D=0
M1789 693 117 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=20370 $D=0
M1790 774 688 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=15740 $D=0
M1791 775 689 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=20370 $D=0
M1792 694 692 774 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=15740 $D=0
M1793 695 693 775 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=20370 $D=0
M1794 167 694 121 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=15740 $D=0
M1795 168 695 122 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=20370 $D=0
M1796 776 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=15740 $D=0
M1797 777 122 168 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=20370 $D=0
M1798 694 690 776 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=15740 $D=0
M1799 695 691 777 168 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=20370 $D=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6 7 8 9 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174
** N=1103 EP=172 IP=2241 FDC=2700
M0 177 1 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 178 1 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=5230 $D=1
M2 179 1 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=9860 $D=1
M3 180 177 2 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=600 $D=1
M4 181 178 3 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=5230 $D=1
M5 182 179 4 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=1045 $Y=9860 $D=1
M6 7 1 180 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=600 $D=1
M7 8 1 181 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=5230 $D=1
M8 9 1 182 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=1565 $Y=9860 $D=1
M9 183 177 5 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=600 $D=1
M10 184 178 5 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=5230 $D=1
M11 185 179 5 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=2375 $Y=9860 $D=1
M12 6 1 183 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=600 $D=1
M13 6 1 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=5230 $D=1
M14 6 1 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=2895 $Y=9860 $D=1
M15 186 177 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=600 $D=1
M16 187 178 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=5230 $D=1
M17 188 179 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3705 $Y=9860 $D=1
M18 7 1 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=600 $D=1
M19 8 1 187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=5230 $D=1
M20 9 1 188 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4225 $Y=9860 $D=1
M21 192 189 186 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=600 $D=1
M22 193 190 187 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=5230 $D=1
M23 194 191 188 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=5035 $Y=9860 $D=1
M24 189 11 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=600 $D=1
M25 190 11 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=5230 $D=1
M26 191 11 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5770 $Y=9860 $D=1
M27 195 189 183 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=600 $D=1
M28 196 190 184 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=5230 $D=1
M29 197 191 185 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=6505 $Y=9860 $D=1
M30 180 11 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=600 $D=1
M31 181 11 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=5230 $D=1
M32 182 11 197 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=7025 $Y=9860 $D=1
M33 198 12 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=600 $D=1
M34 199 12 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=5230 $D=1
M35 200 12 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=7760 $Y=9860 $D=1
M36 201 198 195 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=600 $D=1
M37 202 199 196 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=5230 $D=1
M38 203 200 197 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=8495 $Y=9860 $D=1
M39 192 12 201 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=600 $D=1
M40 193 12 202 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=5230 $D=1
M41 194 12 203 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=9015 $Y=9860 $D=1
M42 204 13 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=600 $D=1
M43 205 13 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=5230 $D=1
M44 206 13 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=9750 $Y=9860 $D=1
M45 207 204 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=600 $D=1
M46 208 205 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=5230 $D=1
M47 209 206 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=10485 $Y=9860 $D=1
M48 14 13 207 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=600 $D=1
M49 15 13 208 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=5230 $D=1
M50 16 13 209 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=11005 $Y=9860 $D=1
M51 210 204 17 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=600 $D=1
M52 211 205 18 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=5230 $D=1
M53 212 206 19 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=11815 $Y=9860 $D=1
M54 213 13 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=600 $D=1
M55 214 13 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=5230 $D=1
M56 215 13 212 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=12335 $Y=9860 $D=1
M57 219 204 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=600 $D=1
M58 220 205 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=5230 $D=1
M59 221 206 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=13145 $Y=9860 $D=1
M60 201 13 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=600 $D=1
M61 202 13 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=5230 $D=1
M62 203 13 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=13665 $Y=9860 $D=1
M63 225 222 219 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=600 $D=1
M64 226 223 220 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=5230 $D=1
M65 227 224 221 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=14475 $Y=9860 $D=1
M66 222 20 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=600 $D=1
M67 223 20 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=5230 $D=1
M68 224 20 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=15210 $Y=9860 $D=1
M69 228 222 210 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=600 $D=1
M70 229 223 211 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=5230 $D=1
M71 230 224 212 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=15945 $Y=9860 $D=1
M72 207 20 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=600 $D=1
M73 208 20 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=5230 $D=1
M74 209 20 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=16465 $Y=9860 $D=1
M75 231 21 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=600 $D=1
M76 232 21 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=5230 $D=1
M77 233 21 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=17200 $Y=9860 $D=1
M78 234 231 228 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=600 $D=1
M79 235 232 229 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=5230 $D=1
M80 236 233 230 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=17935 $Y=9860 $D=1
M81 225 21 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=600 $D=1
M82 226 21 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=5230 $D=1
M83 227 21 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=18455 $Y=9860 $D=1
M84 7 22 237 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=600 $D=1
M85 8 22 238 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=5230 $D=1
M86 9 22 239 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=19190 $Y=9860 $D=1
M87 240 23 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=600 $D=1
M88 241 23 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=5230 $D=1
M89 242 23 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=19570 $Y=9860 $D=1
M90 243 22 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=600 $D=1
M91 244 22 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=5230 $D=1
M92 245 22 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=20305 $Y=9860 $D=1
M93 7 243 951 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=600 $D=1
M94 8 244 952 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=5230 $D=1
M95 9 245 953 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=21040 $Y=9860 $D=1
M96 246 951 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=600 $D=1
M97 247 952 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=5230 $D=1
M98 248 953 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=21420 $Y=9860 $D=1
M99 243 237 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=600 $D=1
M100 244 238 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=5230 $D=1
M101 245 239 248 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=21865 $Y=9860 $D=1
M102 246 23 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=600 $D=1
M103 247 23 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=5230 $D=1
M104 248 23 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=22675 $Y=9860 $D=1
M105 255 24 246 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=600 $D=1
M106 256 24 247 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=5230 $D=1
M107 257 24 248 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=23195 $Y=9860 $D=1
M108 252 24 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=600 $D=1
M109 253 24 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=5230 $D=1
M110 254 24 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=23930 $Y=9860 $D=1
M111 7 25 258 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=600 $D=1
M112 8 25 259 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=5230 $D=1
M113 9 25 260 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=24590 $Y=9860 $D=1
M114 261 26 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=600 $D=1
M115 262 26 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=5230 $D=1
M116 263 26 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=24970 $Y=9860 $D=1
M117 264 25 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=600 $D=1
M118 265 25 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=5230 $D=1
M119 266 25 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=25705 $Y=9860 $D=1
M120 7 264 954 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=600 $D=1
M121 8 265 955 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=5230 $D=1
M122 9 266 956 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=26440 $Y=9860 $D=1
M123 267 954 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=600 $D=1
M124 268 955 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=5230 $D=1
M125 269 956 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=26820 $Y=9860 $D=1
M126 264 258 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=600 $D=1
M127 265 259 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=5230 $D=1
M128 266 260 269 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=27265 $Y=9860 $D=1
M129 267 26 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=600 $D=1
M130 268 26 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=5230 $D=1
M131 269 26 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=28075 $Y=9860 $D=1
M132 255 27 267 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=600 $D=1
M133 256 27 268 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=5230 $D=1
M134 257 27 269 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=28595 $Y=9860 $D=1
M135 270 27 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=600 $D=1
M136 271 27 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=5230 $D=1
M137 272 27 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=29330 $Y=9860 $D=1
M138 7 28 273 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=600 $D=1
M139 8 28 274 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=5230 $D=1
M140 9 28 275 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=29990 $Y=9860 $D=1
M141 276 29 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=600 $D=1
M142 277 29 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=5230 $D=1
M143 278 29 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=30370 $Y=9860 $D=1
M144 279 28 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=600 $D=1
M145 280 28 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=5230 $D=1
M146 281 28 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=31105 $Y=9860 $D=1
M147 7 279 957 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=600 $D=1
M148 8 280 958 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=5230 $D=1
M149 9 281 959 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=31840 $Y=9860 $D=1
M150 282 957 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=600 $D=1
M151 283 958 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=5230 $D=1
M152 284 959 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=32220 $Y=9860 $D=1
M153 279 273 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=600 $D=1
M154 280 274 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=5230 $D=1
M155 281 275 284 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=32665 $Y=9860 $D=1
M156 282 29 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=600 $D=1
M157 283 29 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=5230 $D=1
M158 284 29 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=33475 $Y=9860 $D=1
M159 255 30 282 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=600 $D=1
M160 256 30 283 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=5230 $D=1
M161 257 30 284 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=33995 $Y=9860 $D=1
M162 285 30 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=600 $D=1
M163 286 30 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=5230 $D=1
M164 287 30 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=34730 $Y=9860 $D=1
M165 7 31 288 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=600 $D=1
M166 8 31 289 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=5230 $D=1
M167 9 31 290 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=35390 $Y=9860 $D=1
M168 291 32 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=600 $D=1
M169 292 32 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=5230 $D=1
M170 293 32 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=35770 $Y=9860 $D=1
M171 294 31 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=600 $D=1
M172 295 31 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=5230 $D=1
M173 296 31 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=36505 $Y=9860 $D=1
M174 7 294 960 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=600 $D=1
M175 8 295 961 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=5230 $D=1
M176 9 296 962 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=37240 $Y=9860 $D=1
M177 297 960 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=600 $D=1
M178 298 961 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=5230 $D=1
M179 299 962 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=37620 $Y=9860 $D=1
M180 294 288 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=600 $D=1
M181 295 289 298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=5230 $D=1
M182 296 290 299 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=38065 $Y=9860 $D=1
M183 297 32 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=600 $D=1
M184 298 32 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=5230 $D=1
M185 299 32 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=38875 $Y=9860 $D=1
M186 255 33 297 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=600 $D=1
M187 256 33 298 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=5230 $D=1
M188 257 33 299 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=39395 $Y=9860 $D=1
M189 300 33 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=600 $D=1
M190 301 33 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=5230 $D=1
M191 302 33 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=40130 $Y=9860 $D=1
M192 7 34 303 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=600 $D=1
M193 8 34 304 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=5230 $D=1
M194 9 34 305 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=40790 $Y=9860 $D=1
M195 306 35 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=600 $D=1
M196 307 35 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=5230 $D=1
M197 308 35 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=41170 $Y=9860 $D=1
M198 309 34 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=600 $D=1
M199 310 34 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=5230 $D=1
M200 311 34 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=41905 $Y=9860 $D=1
M201 7 309 963 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=600 $D=1
M202 8 310 964 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=5230 $D=1
M203 9 311 965 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=42640 $Y=9860 $D=1
M204 312 963 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=600 $D=1
M205 313 964 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=5230 $D=1
M206 314 965 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=43020 $Y=9860 $D=1
M207 309 303 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=600 $D=1
M208 310 304 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=5230 $D=1
M209 311 305 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=43465 $Y=9860 $D=1
M210 312 35 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=600 $D=1
M211 313 35 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=5230 $D=1
M212 314 35 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=44275 $Y=9860 $D=1
M213 255 36 312 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=600 $D=1
M214 256 36 313 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=5230 $D=1
M215 257 36 314 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=44795 $Y=9860 $D=1
M216 315 36 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=600 $D=1
M217 316 36 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=5230 $D=1
M218 317 36 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=45530 $Y=9860 $D=1
M219 7 37 318 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=600 $D=1
M220 8 37 319 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=5230 $D=1
M221 9 37 320 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=46190 $Y=9860 $D=1
M222 321 38 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=600 $D=1
M223 322 38 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=5230 $D=1
M224 323 38 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=46570 $Y=9860 $D=1
M225 324 37 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=600 $D=1
M226 325 37 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=5230 $D=1
M227 326 37 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=47305 $Y=9860 $D=1
M228 7 324 966 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=600 $D=1
M229 8 325 967 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=5230 $D=1
M230 9 326 968 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=48040 $Y=9860 $D=1
M231 327 966 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=600 $D=1
M232 328 967 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=5230 $D=1
M233 329 968 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=48420 $Y=9860 $D=1
M234 324 318 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=600 $D=1
M235 325 319 328 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=5230 $D=1
M236 326 320 329 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=48865 $Y=9860 $D=1
M237 327 38 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=600 $D=1
M238 328 38 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=5230 $D=1
M239 329 38 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=49675 $Y=9860 $D=1
M240 255 39 327 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=600 $D=1
M241 256 39 328 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=5230 $D=1
M242 257 39 329 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=50195 $Y=9860 $D=1
M243 330 39 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=600 $D=1
M244 331 39 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=5230 $D=1
M245 332 39 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=50930 $Y=9860 $D=1
M246 7 40 333 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=600 $D=1
M247 8 40 334 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=5230 $D=1
M248 9 40 335 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=51590 $Y=9860 $D=1
M249 336 41 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=600 $D=1
M250 337 41 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=5230 $D=1
M251 338 41 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=51970 $Y=9860 $D=1
M252 339 40 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=600 $D=1
M253 340 40 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=5230 $D=1
M254 341 40 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=52705 $Y=9860 $D=1
M255 7 339 969 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=600 $D=1
M256 8 340 970 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=5230 $D=1
M257 9 341 971 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=53440 $Y=9860 $D=1
M258 342 969 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=600 $D=1
M259 343 970 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=5230 $D=1
M260 344 971 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=53820 $Y=9860 $D=1
M261 339 333 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=600 $D=1
M262 340 334 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=5230 $D=1
M263 341 335 344 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=54265 $Y=9860 $D=1
M264 342 41 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=600 $D=1
M265 343 41 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=5230 $D=1
M266 344 41 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=55075 $Y=9860 $D=1
M267 255 42 342 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=600 $D=1
M268 256 42 343 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=5230 $D=1
M269 257 42 344 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=55595 $Y=9860 $D=1
M270 345 42 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=600 $D=1
M271 346 42 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=5230 $D=1
M272 347 42 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=56330 $Y=9860 $D=1
M273 7 43 348 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=600 $D=1
M274 8 43 349 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=5230 $D=1
M275 9 43 350 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=56990 $Y=9860 $D=1
M276 351 44 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=600 $D=1
M277 352 44 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=5230 $D=1
M278 353 44 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=57370 $Y=9860 $D=1
M279 354 43 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=600 $D=1
M280 355 43 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=5230 $D=1
M281 356 43 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=58105 $Y=9860 $D=1
M282 7 354 972 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=600 $D=1
M283 8 355 973 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=5230 $D=1
M284 9 356 974 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=58840 $Y=9860 $D=1
M285 357 972 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=600 $D=1
M286 358 973 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=5230 $D=1
M287 359 974 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=59220 $Y=9860 $D=1
M288 354 348 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=600 $D=1
M289 355 349 358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=5230 $D=1
M290 356 350 359 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=59665 $Y=9860 $D=1
M291 357 44 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=600 $D=1
M292 358 44 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=5230 $D=1
M293 359 44 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=60475 $Y=9860 $D=1
M294 255 45 357 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=600 $D=1
M295 256 45 358 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=5230 $D=1
M296 257 45 359 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=60995 $Y=9860 $D=1
M297 360 45 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=600 $D=1
M298 361 45 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=5230 $D=1
M299 362 45 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=61730 $Y=9860 $D=1
M300 7 46 363 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=600 $D=1
M301 8 46 364 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=5230 $D=1
M302 9 46 365 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=62390 $Y=9860 $D=1
M303 366 47 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=600 $D=1
M304 367 47 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=5230 $D=1
M305 368 47 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=62770 $Y=9860 $D=1
M306 369 46 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=600 $D=1
M307 370 46 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=5230 $D=1
M308 371 46 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=63505 $Y=9860 $D=1
M309 7 369 975 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=600 $D=1
M310 8 370 976 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=5230 $D=1
M311 9 371 977 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=64240 $Y=9860 $D=1
M312 372 975 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=600 $D=1
M313 373 976 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=5230 $D=1
M314 374 977 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=64620 $Y=9860 $D=1
M315 369 363 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=600 $D=1
M316 370 364 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=5230 $D=1
M317 371 365 374 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=65065 $Y=9860 $D=1
M318 372 47 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=600 $D=1
M319 373 47 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=5230 $D=1
M320 374 47 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=65875 $Y=9860 $D=1
M321 255 48 372 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=600 $D=1
M322 256 48 373 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=5230 $D=1
M323 257 48 374 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=66395 $Y=9860 $D=1
M324 375 48 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=600 $D=1
M325 376 48 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=5230 $D=1
M326 377 48 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=67130 $Y=9860 $D=1
M327 7 49 378 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=600 $D=1
M328 8 49 379 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=5230 $D=1
M329 9 49 380 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=67790 $Y=9860 $D=1
M330 381 50 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=600 $D=1
M331 382 50 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=5230 $D=1
M332 383 50 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=68170 $Y=9860 $D=1
M333 384 49 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=600 $D=1
M334 385 49 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=5230 $D=1
M335 386 49 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=68905 $Y=9860 $D=1
M336 7 384 978 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=600 $D=1
M337 8 385 979 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=5230 $D=1
M338 9 386 980 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=69640 $Y=9860 $D=1
M339 387 978 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=600 $D=1
M340 388 979 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=5230 $D=1
M341 389 980 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=70020 $Y=9860 $D=1
M342 384 378 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=600 $D=1
M343 385 379 388 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=5230 $D=1
M344 386 380 389 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=70465 $Y=9860 $D=1
M345 387 50 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=600 $D=1
M346 388 50 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=5230 $D=1
M347 389 50 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=71275 $Y=9860 $D=1
M348 255 51 387 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=600 $D=1
M349 256 51 388 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=5230 $D=1
M350 257 51 389 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=71795 $Y=9860 $D=1
M351 390 51 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=600 $D=1
M352 391 51 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=5230 $D=1
M353 392 51 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=72530 $Y=9860 $D=1
M354 7 52 393 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=600 $D=1
M355 8 52 394 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=5230 $D=1
M356 9 52 395 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=73190 $Y=9860 $D=1
M357 396 53 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=600 $D=1
M358 397 53 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=5230 $D=1
M359 398 53 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=73570 $Y=9860 $D=1
M360 399 52 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=600 $D=1
M361 400 52 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=5230 $D=1
M362 401 52 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=74305 $Y=9860 $D=1
M363 7 399 981 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=600 $D=1
M364 8 400 982 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=5230 $D=1
M365 9 401 983 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=75040 $Y=9860 $D=1
M366 402 981 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=600 $D=1
M367 403 982 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=5230 $D=1
M368 404 983 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=75420 $Y=9860 $D=1
M369 399 393 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=600 $D=1
M370 400 394 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=5230 $D=1
M371 401 395 404 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=75865 $Y=9860 $D=1
M372 402 53 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=600 $D=1
M373 403 53 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=5230 $D=1
M374 404 53 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=76675 $Y=9860 $D=1
M375 255 54 402 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=600 $D=1
M376 256 54 403 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=5230 $D=1
M377 257 54 404 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=77195 $Y=9860 $D=1
M378 405 54 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=600 $D=1
M379 406 54 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=5230 $D=1
M380 407 54 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=77930 $Y=9860 $D=1
M381 7 55 408 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=600 $D=1
M382 8 55 409 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=5230 $D=1
M383 9 55 410 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=78590 $Y=9860 $D=1
M384 411 56 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=600 $D=1
M385 412 56 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=5230 $D=1
M386 413 56 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=78970 $Y=9860 $D=1
M387 414 55 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=600 $D=1
M388 415 55 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=5230 $D=1
M389 416 55 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=79705 $Y=9860 $D=1
M390 7 414 984 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=600 $D=1
M391 8 415 985 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=5230 $D=1
M392 9 416 986 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=80440 $Y=9860 $D=1
M393 417 984 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=600 $D=1
M394 418 985 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=5230 $D=1
M395 419 986 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=80820 $Y=9860 $D=1
M396 414 408 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=600 $D=1
M397 415 409 418 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=5230 $D=1
M398 416 410 419 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=81265 $Y=9860 $D=1
M399 417 56 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=600 $D=1
M400 418 56 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=5230 $D=1
M401 419 56 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=82075 $Y=9860 $D=1
M402 255 57 417 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=600 $D=1
M403 256 57 418 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=5230 $D=1
M404 257 57 419 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=82595 $Y=9860 $D=1
M405 420 57 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=600 $D=1
M406 421 57 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=5230 $D=1
M407 422 57 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=83330 $Y=9860 $D=1
M408 7 58 423 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=600 $D=1
M409 8 58 424 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=5230 $D=1
M410 9 58 425 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=83990 $Y=9860 $D=1
M411 426 59 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=600 $D=1
M412 427 59 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=5230 $D=1
M413 428 59 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=84370 $Y=9860 $D=1
M414 429 58 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=600 $D=1
M415 430 58 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=5230 $D=1
M416 431 58 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=85105 $Y=9860 $D=1
M417 7 429 987 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=600 $D=1
M418 8 430 988 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=5230 $D=1
M419 9 431 989 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=85840 $Y=9860 $D=1
M420 432 987 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=600 $D=1
M421 433 988 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=5230 $D=1
M422 434 989 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=86220 $Y=9860 $D=1
M423 429 423 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=600 $D=1
M424 430 424 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=5230 $D=1
M425 431 425 434 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=86665 $Y=9860 $D=1
M426 432 59 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=600 $D=1
M427 433 59 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=5230 $D=1
M428 434 59 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=87475 $Y=9860 $D=1
M429 255 60 432 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=600 $D=1
M430 256 60 433 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=5230 $D=1
M431 257 60 434 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=87995 $Y=9860 $D=1
M432 435 60 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=600 $D=1
M433 436 60 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=5230 $D=1
M434 437 60 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=88730 $Y=9860 $D=1
M435 7 61 438 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=600 $D=1
M436 8 61 439 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=5230 $D=1
M437 9 61 440 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=89390 $Y=9860 $D=1
M438 441 62 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=600 $D=1
M439 442 62 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=5230 $D=1
M440 443 62 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=89770 $Y=9860 $D=1
M441 444 61 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=600 $D=1
M442 445 61 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=5230 $D=1
M443 446 61 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=90505 $Y=9860 $D=1
M444 7 444 990 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=600 $D=1
M445 8 445 991 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=5230 $D=1
M446 9 446 992 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=91240 $Y=9860 $D=1
M447 447 990 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=600 $D=1
M448 448 991 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=5230 $D=1
M449 449 992 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=91620 $Y=9860 $D=1
M450 444 438 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=600 $D=1
M451 445 439 448 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=5230 $D=1
M452 446 440 449 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=92065 $Y=9860 $D=1
M453 447 62 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=600 $D=1
M454 448 62 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=5230 $D=1
M455 449 62 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=92875 $Y=9860 $D=1
M456 255 63 447 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=600 $D=1
M457 256 63 448 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=5230 $D=1
M458 257 63 449 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=93395 $Y=9860 $D=1
M459 450 63 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=600 $D=1
M460 451 63 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=5230 $D=1
M461 452 63 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=94130 $Y=9860 $D=1
M462 7 64 453 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=600 $D=1
M463 8 64 454 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=5230 $D=1
M464 9 64 455 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=94790 $Y=9860 $D=1
M465 456 65 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=600 $D=1
M466 457 65 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=5230 $D=1
M467 458 65 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=95170 $Y=9860 $D=1
M468 459 64 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=600 $D=1
M469 460 64 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=5230 $D=1
M470 461 64 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=95905 $Y=9860 $D=1
M471 7 459 993 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=600 $D=1
M472 8 460 994 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=5230 $D=1
M473 9 461 995 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=96640 $Y=9860 $D=1
M474 462 993 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=600 $D=1
M475 463 994 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=5230 $D=1
M476 464 995 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=97020 $Y=9860 $D=1
M477 459 453 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=600 $D=1
M478 460 454 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=5230 $D=1
M479 461 455 464 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=97465 $Y=9860 $D=1
M480 462 65 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=600 $D=1
M481 463 65 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=5230 $D=1
M482 464 65 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=98275 $Y=9860 $D=1
M483 255 66 462 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=600 $D=1
M484 256 66 463 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=5230 $D=1
M485 257 66 464 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=98795 $Y=9860 $D=1
M486 465 66 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=600 $D=1
M487 466 66 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=5230 $D=1
M488 467 66 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=99530 $Y=9860 $D=1
M489 7 67 468 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=600 $D=1
M490 8 67 469 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=5230 $D=1
M491 9 67 470 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=100190 $Y=9860 $D=1
M492 471 68 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=600 $D=1
M493 472 68 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=5230 $D=1
M494 473 68 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=100570 $Y=9860 $D=1
M495 474 67 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=600 $D=1
M496 475 67 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=5230 $D=1
M497 476 67 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=101305 $Y=9860 $D=1
M498 7 474 996 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=600 $D=1
M499 8 475 997 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=5230 $D=1
M500 9 476 998 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=102040 $Y=9860 $D=1
M501 477 996 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=600 $D=1
M502 478 997 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=5230 $D=1
M503 479 998 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=102420 $Y=9860 $D=1
M504 474 468 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=600 $D=1
M505 475 469 478 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=5230 $D=1
M506 476 470 479 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=102865 $Y=9860 $D=1
M507 477 68 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=600 $D=1
M508 478 68 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=5230 $D=1
M509 479 68 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=103675 $Y=9860 $D=1
M510 255 69 477 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=600 $D=1
M511 256 69 478 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=5230 $D=1
M512 257 69 479 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=104195 $Y=9860 $D=1
M513 480 69 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=600 $D=1
M514 481 69 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=5230 $D=1
M515 482 69 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=104930 $Y=9860 $D=1
M516 7 70 483 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=600 $D=1
M517 8 70 484 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=5230 $D=1
M518 9 70 485 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=105590 $Y=9860 $D=1
M519 486 71 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=600 $D=1
M520 487 71 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=5230 $D=1
M521 488 71 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=105970 $Y=9860 $D=1
M522 489 70 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=600 $D=1
M523 490 70 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=5230 $D=1
M524 491 70 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=106705 $Y=9860 $D=1
M525 7 489 999 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=600 $D=1
M526 8 490 1000 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=5230 $D=1
M527 9 491 1001 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=107440 $Y=9860 $D=1
M528 492 999 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=600 $D=1
M529 493 1000 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=5230 $D=1
M530 494 1001 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=107820 $Y=9860 $D=1
M531 489 483 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=600 $D=1
M532 490 484 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=5230 $D=1
M533 491 485 494 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=108265 $Y=9860 $D=1
M534 492 71 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=600 $D=1
M535 493 71 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=5230 $D=1
M536 494 71 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=109075 $Y=9860 $D=1
M537 255 72 492 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=600 $D=1
M538 256 72 493 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=5230 $D=1
M539 257 72 494 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=109595 $Y=9860 $D=1
M540 495 72 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=600 $D=1
M541 496 72 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=5230 $D=1
M542 497 72 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=110330 $Y=9860 $D=1
M543 7 73 498 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=600 $D=1
M544 8 73 499 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=5230 $D=1
M545 9 73 500 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=110990 $Y=9860 $D=1
M546 501 74 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=600 $D=1
M547 502 74 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=5230 $D=1
M548 503 74 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=111370 $Y=9860 $D=1
M549 504 73 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=600 $D=1
M550 505 73 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=5230 $D=1
M551 506 73 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=112105 $Y=9860 $D=1
M552 7 504 1002 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=600 $D=1
M553 8 505 1003 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=5230 $D=1
M554 9 506 1004 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=112840 $Y=9860 $D=1
M555 507 1002 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=600 $D=1
M556 508 1003 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=5230 $D=1
M557 509 1004 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=113220 $Y=9860 $D=1
M558 504 498 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=600 $D=1
M559 505 499 508 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=5230 $D=1
M560 506 500 509 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=113665 $Y=9860 $D=1
M561 507 74 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=600 $D=1
M562 508 74 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=5230 $D=1
M563 509 74 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=114475 $Y=9860 $D=1
M564 255 75 507 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=600 $D=1
M565 256 75 508 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=5230 $D=1
M566 257 75 509 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=114995 $Y=9860 $D=1
M567 510 75 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=600 $D=1
M568 511 75 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=5230 $D=1
M569 512 75 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=115730 $Y=9860 $D=1
M570 7 76 513 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=600 $D=1
M571 8 76 514 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=5230 $D=1
M572 9 76 515 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=116390 $Y=9860 $D=1
M573 516 77 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=600 $D=1
M574 517 77 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=5230 $D=1
M575 518 77 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=116770 $Y=9860 $D=1
M576 519 76 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=600 $D=1
M577 520 76 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=5230 $D=1
M578 521 76 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=117505 $Y=9860 $D=1
M579 7 519 1005 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=600 $D=1
M580 8 520 1006 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=5230 $D=1
M581 9 521 1007 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=118240 $Y=9860 $D=1
M582 522 1005 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=600 $D=1
M583 523 1006 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=5230 $D=1
M584 524 1007 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=118620 $Y=9860 $D=1
M585 519 513 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=600 $D=1
M586 520 514 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=5230 $D=1
M587 521 515 524 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=119065 $Y=9860 $D=1
M588 522 77 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=600 $D=1
M589 523 77 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=5230 $D=1
M590 524 77 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=119875 $Y=9860 $D=1
M591 255 78 522 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=600 $D=1
M592 256 78 523 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=5230 $D=1
M593 257 78 524 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=120395 $Y=9860 $D=1
M594 525 78 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=600 $D=1
M595 526 78 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=5230 $D=1
M596 527 78 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=121130 $Y=9860 $D=1
M597 7 79 528 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=600 $D=1
M598 8 79 529 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=5230 $D=1
M599 9 79 530 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=121790 $Y=9860 $D=1
M600 531 80 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=600 $D=1
M601 532 80 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=5230 $D=1
M602 533 80 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=122170 $Y=9860 $D=1
M603 534 79 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=600 $D=1
M604 535 79 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=5230 $D=1
M605 536 79 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=122905 $Y=9860 $D=1
M606 7 534 1008 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=600 $D=1
M607 8 535 1009 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=5230 $D=1
M608 9 536 1010 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=123640 $Y=9860 $D=1
M609 537 1008 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=600 $D=1
M610 538 1009 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=5230 $D=1
M611 539 1010 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=124020 $Y=9860 $D=1
M612 534 528 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=600 $D=1
M613 535 529 538 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=5230 $D=1
M614 536 530 539 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=124465 $Y=9860 $D=1
M615 537 80 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=600 $D=1
M616 538 80 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=5230 $D=1
M617 539 80 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=125275 $Y=9860 $D=1
M618 255 81 537 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=600 $D=1
M619 256 81 538 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=5230 $D=1
M620 257 81 539 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=125795 $Y=9860 $D=1
M621 540 81 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=600 $D=1
M622 541 81 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=5230 $D=1
M623 542 81 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=126530 $Y=9860 $D=1
M624 7 82 543 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=600 $D=1
M625 8 82 544 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=5230 $D=1
M626 9 82 545 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=127190 $Y=9860 $D=1
M627 546 83 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=600 $D=1
M628 547 83 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=5230 $D=1
M629 548 83 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=127570 $Y=9860 $D=1
M630 549 82 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=600 $D=1
M631 550 82 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=5230 $D=1
M632 551 82 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=128305 $Y=9860 $D=1
M633 7 549 1011 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=600 $D=1
M634 8 550 1012 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=5230 $D=1
M635 9 551 1013 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=129040 $Y=9860 $D=1
M636 552 1011 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=600 $D=1
M637 553 1012 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=5230 $D=1
M638 554 1013 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=129420 $Y=9860 $D=1
M639 549 543 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=600 $D=1
M640 550 544 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=5230 $D=1
M641 551 545 554 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=129865 $Y=9860 $D=1
M642 552 83 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=600 $D=1
M643 553 83 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=5230 $D=1
M644 554 83 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=130675 $Y=9860 $D=1
M645 255 84 552 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=600 $D=1
M646 256 84 553 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=5230 $D=1
M647 257 84 554 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=131195 $Y=9860 $D=1
M648 555 84 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=600 $D=1
M649 556 84 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=5230 $D=1
M650 557 84 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=131930 $Y=9860 $D=1
M651 7 85 558 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=600 $D=1
M652 8 85 559 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=5230 $D=1
M653 9 85 560 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=132590 $Y=9860 $D=1
M654 561 86 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=600 $D=1
M655 562 86 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=5230 $D=1
M656 563 86 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=132970 $Y=9860 $D=1
M657 564 85 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=600 $D=1
M658 565 85 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=5230 $D=1
M659 566 85 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=133705 $Y=9860 $D=1
M660 7 564 1014 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=600 $D=1
M661 8 565 1015 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=5230 $D=1
M662 9 566 1016 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=134440 $Y=9860 $D=1
M663 567 1014 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=600 $D=1
M664 568 1015 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=5230 $D=1
M665 569 1016 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=134820 $Y=9860 $D=1
M666 564 558 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=600 $D=1
M667 565 559 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=5230 $D=1
M668 566 560 569 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=135265 $Y=9860 $D=1
M669 567 86 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=600 $D=1
M670 568 86 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=5230 $D=1
M671 569 86 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=136075 $Y=9860 $D=1
M672 255 87 567 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=600 $D=1
M673 256 87 568 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=5230 $D=1
M674 257 87 569 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=136595 $Y=9860 $D=1
M675 570 87 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=600 $D=1
M676 571 87 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=5230 $D=1
M677 572 87 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=137330 $Y=9860 $D=1
M678 7 88 573 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=600 $D=1
M679 8 88 574 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=5230 $D=1
M680 9 88 575 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=137990 $Y=9860 $D=1
M681 576 89 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=600 $D=1
M682 577 89 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=5230 $D=1
M683 578 89 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=138370 $Y=9860 $D=1
M684 579 88 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=600 $D=1
M685 580 88 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=5230 $D=1
M686 581 88 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=139105 $Y=9860 $D=1
M687 7 579 1017 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=600 $D=1
M688 8 580 1018 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=5230 $D=1
M689 9 581 1019 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=139840 $Y=9860 $D=1
M690 582 1017 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=600 $D=1
M691 583 1018 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=5230 $D=1
M692 584 1019 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=140220 $Y=9860 $D=1
M693 579 573 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=600 $D=1
M694 580 574 583 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=5230 $D=1
M695 581 575 584 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=140665 $Y=9860 $D=1
M696 582 89 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=600 $D=1
M697 583 89 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=5230 $D=1
M698 584 89 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=141475 $Y=9860 $D=1
M699 255 90 582 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=600 $D=1
M700 256 90 583 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=5230 $D=1
M701 257 90 584 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=141995 $Y=9860 $D=1
M702 585 90 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=600 $D=1
M703 586 90 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=5230 $D=1
M704 587 90 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=142730 $Y=9860 $D=1
M705 7 91 588 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=600 $D=1
M706 8 91 589 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=5230 $D=1
M707 9 91 590 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=143390 $Y=9860 $D=1
M708 591 92 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=600 $D=1
M709 592 92 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=5230 $D=1
M710 593 92 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=143770 $Y=9860 $D=1
M711 594 91 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=600 $D=1
M712 595 91 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=5230 $D=1
M713 596 91 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=144505 $Y=9860 $D=1
M714 7 594 1020 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=600 $D=1
M715 8 595 1021 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=5230 $D=1
M716 9 596 1022 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=145240 $Y=9860 $D=1
M717 597 1020 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=600 $D=1
M718 598 1021 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=5230 $D=1
M719 599 1022 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=145620 $Y=9860 $D=1
M720 594 588 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=600 $D=1
M721 595 589 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=5230 $D=1
M722 596 590 599 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=146065 $Y=9860 $D=1
M723 597 92 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=600 $D=1
M724 598 92 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=5230 $D=1
M725 599 92 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=146875 $Y=9860 $D=1
M726 255 93 597 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=600 $D=1
M727 256 93 598 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=5230 $D=1
M728 257 93 599 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=147395 $Y=9860 $D=1
M729 600 93 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=600 $D=1
M730 601 93 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=5230 $D=1
M731 602 93 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=148130 $Y=9860 $D=1
M732 7 94 603 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=600 $D=1
M733 8 94 604 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=5230 $D=1
M734 9 94 605 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=148790 $Y=9860 $D=1
M735 606 95 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=600 $D=1
M736 607 95 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=5230 $D=1
M737 608 95 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=149170 $Y=9860 $D=1
M738 609 94 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=600 $D=1
M739 610 94 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=5230 $D=1
M740 611 94 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=149905 $Y=9860 $D=1
M741 7 609 1023 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=600 $D=1
M742 8 610 1024 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=5230 $D=1
M743 9 611 1025 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=150640 $Y=9860 $D=1
M744 612 1023 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=600 $D=1
M745 613 1024 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=5230 $D=1
M746 614 1025 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=151020 $Y=9860 $D=1
M747 609 603 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=600 $D=1
M748 610 604 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=5230 $D=1
M749 611 605 614 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=151465 $Y=9860 $D=1
M750 612 95 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=600 $D=1
M751 613 95 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=5230 $D=1
M752 614 95 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=152275 $Y=9860 $D=1
M753 255 96 612 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=600 $D=1
M754 256 96 613 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=5230 $D=1
M755 257 96 614 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=152795 $Y=9860 $D=1
M756 615 96 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=600 $D=1
M757 616 96 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=5230 $D=1
M758 617 96 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=153530 $Y=9860 $D=1
M759 7 97 618 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=600 $D=1
M760 8 97 619 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=5230 $D=1
M761 9 97 620 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=154190 $Y=9860 $D=1
M762 621 98 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=600 $D=1
M763 622 98 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=5230 $D=1
M764 623 98 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=154570 $Y=9860 $D=1
M765 624 97 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=600 $D=1
M766 625 97 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=5230 $D=1
M767 626 97 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=155305 $Y=9860 $D=1
M768 7 624 1026 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=600 $D=1
M769 8 625 1027 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=5230 $D=1
M770 9 626 1028 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=156040 $Y=9860 $D=1
M771 627 1026 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=600 $D=1
M772 628 1027 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=5230 $D=1
M773 629 1028 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=156420 $Y=9860 $D=1
M774 624 618 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=600 $D=1
M775 625 619 628 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=5230 $D=1
M776 626 620 629 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=156865 $Y=9860 $D=1
M777 627 98 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=600 $D=1
M778 628 98 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=5230 $D=1
M779 629 98 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=157675 $Y=9860 $D=1
M780 255 99 627 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=600 $D=1
M781 256 99 628 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=5230 $D=1
M782 257 99 629 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=158195 $Y=9860 $D=1
M783 630 99 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=600 $D=1
M784 631 99 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=5230 $D=1
M785 632 99 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=158930 $Y=9860 $D=1
M786 7 100 633 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=600 $D=1
M787 8 100 634 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=5230 $D=1
M788 9 100 635 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=159590 $Y=9860 $D=1
M789 636 101 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=600 $D=1
M790 637 101 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=5230 $D=1
M791 638 101 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=159970 $Y=9860 $D=1
M792 639 100 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=600 $D=1
M793 640 100 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=5230 $D=1
M794 641 100 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=160705 $Y=9860 $D=1
M795 7 639 1029 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=600 $D=1
M796 8 640 1030 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=5230 $D=1
M797 9 641 1031 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=161440 $Y=9860 $D=1
M798 642 1029 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=600 $D=1
M799 643 1030 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=5230 $D=1
M800 644 1031 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=161820 $Y=9860 $D=1
M801 639 633 642 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=600 $D=1
M802 640 634 643 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=5230 $D=1
M803 641 635 644 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=162265 $Y=9860 $D=1
M804 642 101 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=600 $D=1
M805 643 101 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=5230 $D=1
M806 644 101 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=163075 $Y=9860 $D=1
M807 255 102 642 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=600 $D=1
M808 256 102 643 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=5230 $D=1
M809 257 102 644 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=163595 $Y=9860 $D=1
M810 645 102 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=600 $D=1
M811 646 102 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=5230 $D=1
M812 647 102 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=164330 $Y=9860 $D=1
M813 7 103 648 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=600 $D=1
M814 8 103 649 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=5230 $D=1
M815 9 103 650 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=164990 $Y=9860 $D=1
M816 651 104 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=600 $D=1
M817 652 104 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=5230 $D=1
M818 653 104 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=165370 $Y=9860 $D=1
M819 654 103 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=600 $D=1
M820 655 103 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=5230 $D=1
M821 656 103 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=166105 $Y=9860 $D=1
M822 7 654 1032 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=600 $D=1
M823 8 655 1033 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=5230 $D=1
M824 9 656 1034 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=166840 $Y=9860 $D=1
M825 657 1032 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=600 $D=1
M826 658 1033 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=5230 $D=1
M827 659 1034 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=167220 $Y=9860 $D=1
M828 654 648 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=600 $D=1
M829 655 649 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=5230 $D=1
M830 656 650 659 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=167665 $Y=9860 $D=1
M831 657 104 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=600 $D=1
M832 658 104 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=5230 $D=1
M833 659 104 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=168475 $Y=9860 $D=1
M834 255 105 657 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=600 $D=1
M835 256 105 658 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=5230 $D=1
M836 257 105 659 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=168995 $Y=9860 $D=1
M837 660 105 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=600 $D=1
M838 661 105 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=5230 $D=1
M839 662 105 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=169730 $Y=9860 $D=1
M840 7 106 663 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=600 $D=1
M841 8 106 664 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=5230 $D=1
M842 9 106 665 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=170390 $Y=9860 $D=1
M843 666 107 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=600 $D=1
M844 667 107 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=5230 $D=1
M845 668 107 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=170770 $Y=9860 $D=1
M846 669 106 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=600 $D=1
M847 670 106 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=5230 $D=1
M848 671 106 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=171505 $Y=9860 $D=1
M849 7 669 1035 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=600 $D=1
M850 8 670 1036 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=5230 $D=1
M851 9 671 1037 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=172240 $Y=9860 $D=1
M852 672 1035 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=600 $D=1
M853 673 1036 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=5230 $D=1
M854 674 1037 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=172620 $Y=9860 $D=1
M855 669 663 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=600 $D=1
M856 670 664 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=5230 $D=1
M857 671 665 674 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=173065 $Y=9860 $D=1
M858 672 107 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=600 $D=1
M859 673 107 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=5230 $D=1
M860 674 107 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=173875 $Y=9860 $D=1
M861 255 108 672 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=600 $D=1
M862 256 108 673 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=5230 $D=1
M863 257 108 674 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=174395 $Y=9860 $D=1
M864 675 108 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=600 $D=1
M865 676 108 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=5230 $D=1
M866 677 108 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=175130 $Y=9860 $D=1
M867 7 109 678 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=600 $D=1
M868 8 109 679 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=5230 $D=1
M869 9 109 680 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=175790 $Y=9860 $D=1
M870 681 110 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=600 $D=1
M871 682 110 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=5230 $D=1
M872 683 110 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=176170 $Y=9860 $D=1
M873 684 109 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=600 $D=1
M874 685 109 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=5230 $D=1
M875 686 109 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=176905 $Y=9860 $D=1
M876 7 684 1038 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=600 $D=1
M877 8 685 1039 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=5230 $D=1
M878 9 686 1040 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=177640 $Y=9860 $D=1
M879 687 1038 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=600 $D=1
M880 688 1039 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=5230 $D=1
M881 689 1040 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=178020 $Y=9860 $D=1
M882 684 678 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=600 $D=1
M883 685 679 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=5230 $D=1
M884 686 680 689 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=178465 $Y=9860 $D=1
M885 687 110 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=600 $D=1
M886 688 110 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=5230 $D=1
M887 689 110 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=179275 $Y=9860 $D=1
M888 255 113 687 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=600 $D=1
M889 256 113 688 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=5230 $D=1
M890 257 113 689 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=179795 $Y=9860 $D=1
M891 690 113 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=600 $D=1
M892 691 113 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=5230 $D=1
M893 692 113 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=180530 $Y=9860 $D=1
M894 7 114 693 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=600 $D=1
M895 8 114 694 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=5230 $D=1
M896 9 114 695 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=181190 $Y=9860 $D=1
M897 696 115 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=600 $D=1
M898 697 115 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=5230 $D=1
M899 698 115 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=181570 $Y=9860 $D=1
M900 699 114 234 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=600 $D=1
M901 700 114 235 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=5230 $D=1
M902 701 114 236 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=182305 $Y=9860 $D=1
M903 7 699 1041 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=600 $D=1
M904 8 700 1042 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=5230 $D=1
M905 9 701 1043 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=183040 $Y=9860 $D=1
M906 702 1041 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=600 $D=1
M907 703 1042 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=5230 $D=1
M908 704 1043 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=183420 $Y=9860 $D=1
M909 699 693 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=600 $D=1
M910 700 694 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=5230 $D=1
M911 701 695 704 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=183865 $Y=9860 $D=1
M912 702 115 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=600 $D=1
M913 703 115 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=5230 $D=1
M914 704 115 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=184675 $Y=9860 $D=1
M915 255 118 702 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=600 $D=1
M916 256 118 703 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=5230 $D=1
M917 257 118 704 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=185195 $Y=9860 $D=1
M918 705 118 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=600 $D=1
M919 706 118 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=5230 $D=1
M920 707 118 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=185930 $Y=9860 $D=1
M921 7 119 708 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=600 $D=1
M922 8 119 709 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=5230 $D=1
M923 9 119 710 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=186590 $Y=9860 $D=1
M924 711 120 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=600 $D=1
M925 712 120 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=5230 $D=1
M926 713 120 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=186970 $Y=9860 $D=1
M927 7 120 249 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=600 $D=1
M928 8 120 250 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=5230 $D=1
M929 9 120 251 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=187705 $Y=9860 $D=1
M930 255 119 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=600 $D=1
M931 256 119 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=5230 $D=1
M932 257 119 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=188225 $Y=9860 $D=1
M933 7 717 714 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=600 $D=1
M934 8 718 715 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=5230 $D=1
M935 9 719 716 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=188960 $Y=9860 $D=1
M936 717 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=600 $D=1
M937 718 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=5230 $D=1
M938 719 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=189340 $Y=9860 $D=1
M939 1044 249 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=600 $D=1
M940 1045 250 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=5230 $D=1
M941 1046 251 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=190000 $Y=9860 $D=1
M942 720 714 1044 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=600 $D=1
M943 721 715 1045 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=5230 $D=1
M944 722 716 1046 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=190445 $Y=9860 $D=1
M945 7 720 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=600 $D=1
M946 8 721 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=5230 $D=1
M947 9 722 724 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=191180 $Y=9860 $D=1
M948 1047 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=600 $D=1
M949 1048 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=5230 $D=1
M950 1049 724 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=191560 $Y=9860 $D=1
M951 720 717 1047 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=600 $D=1
M952 721 718 1048 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=5230 $D=1
M953 722 719 1049 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=191940 $Y=9860 $D=1
M954 7 728 725 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=600 $D=1
M955 8 729 726 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=5230 $D=1
M956 9 730 727 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=192955 $Y=9860 $D=1
M957 728 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=600 $D=1
M958 729 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=5230 $D=1
M959 730 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=193335 $Y=9860 $D=1
M960 1050 255 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=600 $D=1
M961 1051 256 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=5230 $D=1
M962 1052 257 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=193995 $Y=9860 $D=1
M963 731 725 1050 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=600 $D=1
M964 732 726 1051 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=5230 $D=1
M965 733 727 1052 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=194440 $Y=9860 $D=1
M966 7 731 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=600 $D=1
M967 8 732 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=5230 $D=1
M968 9 733 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=195175 $Y=9860 $D=1
M969 1053 123 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=600 $D=1
M970 1054 124 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=5230 $D=1
M971 1055 125 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=195555 $Y=9860 $D=1
M972 731 728 1053 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=600 $D=1
M973 732 729 1054 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=5230 $D=1
M974 733 730 1055 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=195935 $Y=9860 $D=1
M975 734 126 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=600 $D=1
M976 735 126 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=5230 $D=1
M977 736 126 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=196950 $Y=9860 $D=1
M978 737 734 122 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=600 $D=1
M979 738 735 723 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=5230 $D=1
M980 739 736 724 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=197685 $Y=9860 $D=1
M981 127 126 737 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=600 $D=1
M982 128 126 738 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=5230 $D=1
M983 129 126 739 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=198205 $Y=9860 $D=1
M984 740 130 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=600 $D=1
M985 741 130 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=5230 $D=1
M986 742 130 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=198945 $Y=9860 $D=1
M987 743 740 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=600 $D=1
M988 744 741 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=5230 $D=1
M989 745 742 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=199680 $Y=9860 $D=1
M990 1056 130 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=600 $D=1
M991 1057 130 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=5230 $D=1
M992 1058 130 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.89e-14 PD=5.25e-07 PS=6e-07 $X=200200 $Y=9860 $D=1
M993 7 123 1056 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=600 $D=1
M994 8 124 1057 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=5230 $D=1
M995 9 125 1058 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.5525e-14 PD=3.8e-07 PS=5.25e-07 $X=200645 $Y=9860 $D=1
M996 746 131 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=600 $D=1
M997 747 131 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=5230 $D=1
M998 748 131 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=201305 $Y=9860 $D=1
M999 749 746 743 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=600 $D=1
M1000 750 747 744 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=5230 $D=1
M1001 751 748 745 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=202040 $Y=9860 $D=1
M1002 14 131 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=600 $D=1
M1003 15 131 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=5230 $D=1
M1004 16 131 751 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=202560 $Y=9860 $D=1
M1005 755 752 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=600 $D=1
M1006 756 753 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=5230 $D=1
M1007 757 754 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=203300 $Y=9860 $D=1
M1008 7 761 758 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=600 $D=1
M1009 8 762 759 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=5230 $D=1
M1010 9 763 760 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=203960 $Y=9860 $D=1
M1011 764 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=600 $D=1
M1012 765 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=5230 $D=1
M1013 766 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=204340 $Y=9860 $D=1
M1014 761 764 752 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=600 $D=1
M1015 762 765 753 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=5230 $D=1
M1016 763 766 754 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=205075 $Y=9860 $D=1
M1017 755 737 761 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=600 $D=1
M1018 756 738 762 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=5230 $D=1
M1019 757 739 763 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=205595 $Y=9860 $D=1
M1020 767 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=600 $D=1
M1021 768 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=5230 $D=1
M1022 769 760 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=206330 $Y=9860 $D=1
M1023 770 767 749 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=600 $D=1
M1024 771 768 750 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=5230 $D=1
M1025 772 769 751 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=207065 $Y=9860 $D=1
M1026 737 758 770 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=600 $D=1
M1027 738 759 771 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=5230 $D=1
M1028 739 760 772 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=207585 $Y=9860 $D=1
M1029 773 770 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=600 $D=1
M1030 774 771 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=5230 $D=1
M1031 775 772 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208320 $Y=9860 $D=1
M1032 776 758 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=600 $D=1
M1033 777 759 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=5230 $D=1
M1034 778 760 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=208980 $Y=9860 $D=1
M1035 779 776 773 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=600 $D=1
M1036 780 777 774 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=5230 $D=1
M1037 781 778 775 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=209715 $Y=9860 $D=1
M1038 749 758 779 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=600 $D=1
M1039 750 759 780 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=5230 $D=1
M1040 751 760 781 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=210235 $Y=9860 $D=1
M1041 782 737 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=600 $D=1
M1042 783 738 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=5230 $D=1
M1043 784 739 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=210970 $Y=9860 $D=1
M1044 7 749 782 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=600 $D=1
M1045 8 750 783 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=5230 $D=1
M1046 9 751 784 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=211350 $Y=9860 $D=1
M1047 785 779 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=600 $D=1
M1048 786 780 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=5230 $D=1
M1049 787 781 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=212010 $Y=9860 $D=1
M1050 1086 737 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=600 $D=1
M1051 1087 738 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=5230 $D=1
M1052 1088 739 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=9860 $D=1
M1053 788 749 1086 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=600 $D=1
M1054 789 750 1087 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=5230 $D=1
M1055 790 751 1088 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=9860 $D=1
M1056 1089 737 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=600 $D=1
M1057 1090 738 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=5230 $D=1
M1058 1091 739 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=9860 $D=1
M1059 791 749 1089 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=600 $D=1
M1060 792 750 1090 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=5230 $D=1
M1061 793 751 1091 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=9860 $D=1
M1062 797 737 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=600 $D=1
M1063 798 738 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=5230 $D=1
M1064 799 739 796 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=214750 $Y=9860 $D=1
M1065 794 749 797 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=600 $D=1
M1066 795 750 798 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=5230 $D=1
M1067 796 751 799 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=215130 $Y=9860 $D=1
M1068 7 791 794 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=600 $D=1
M1069 8 792 795 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=5230 $D=1
M1070 9 793 796 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=2.835e-14 PD=5.65e-07 PS=6.75e-07 $X=215545 $Y=9860 $D=1
M1071 800 135 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=600 $D=1
M1072 801 135 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=5230 $D=1
M1073 802 135 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=216210 $Y=9860 $D=1
M1074 803 800 782 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=600 $D=1
M1075 804 801 783 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=5230 $D=1
M1076 805 802 784 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=216945 $Y=9860 $D=1
M1077 788 135 803 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=600 $D=1
M1078 789 135 804 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=5230 $D=1
M1079 790 135 805 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=217465 $Y=9860 $D=1
M1080 806 800 785 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=600 $D=1
M1081 807 801 786 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=5230 $D=1
M1082 808 802 787 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=218275 $Y=9860 $D=1
M1083 797 135 806 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=600 $D=1
M1084 798 135 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=5230 $D=1
M1085 799 135 808 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=218795 $Y=9860 $D=1
M1086 809 136 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=600 $D=1
M1087 810 136 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=5230 $D=1
M1088 811 136 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=219530 $Y=9860 $D=1
M1089 812 809 806 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=600 $D=1
M1090 813 810 807 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=5230 $D=1
M1091 814 811 808 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=220265 $Y=9860 $D=1
M1092 803 136 812 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=600 $D=1
M1093 804 136 813 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=5230 $D=1
M1094 805 136 814 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=220785 $Y=9860 $D=1
M1095 17 812 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=600 $D=1
M1096 18 813 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=5230 $D=1
M1097 19 814 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=221520 $Y=9860 $D=1
M1098 815 137 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=600 $D=1
M1099 816 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=5230 $D=1
M1100 817 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=222180 $Y=9860 $D=1
M1101 818 815 138 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=600 $D=1
M1102 819 816 139 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=5230 $D=1
M1103 820 817 140 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=222915 $Y=9860 $D=1
M1104 141 137 818 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=600 $D=1
M1105 142 137 819 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=5230 $D=1
M1106 138 137 820 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=223435 $Y=9860 $D=1
M1107 821 137 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=600 $D=1
M1108 822 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=5230 $D=1
M1109 823 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=224170 $Y=9860 $D=1
M1110 824 821 143 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=600 $D=1
M1111 825 822 144 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=5230 $D=1
M1112 826 823 145 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=224905 $Y=9860 $D=1
M1113 141 137 824 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=600 $D=1
M1114 141 137 825 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=5230 $D=1
M1115 146 137 826 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=225425 $Y=9860 $D=1
M1116 827 137 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=600 $D=1
M1117 828 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=5230 $D=1
M1118 829 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=226160 $Y=9860 $D=1
M1119 830 827 134 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=600 $D=1
M1120 831 828 133 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=5230 $D=1
M1121 832 829 132 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=226895 $Y=9860 $D=1
M1122 141 137 830 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=600 $D=1
M1123 141 137 831 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=5230 $D=1
M1124 141 137 832 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=227415 $Y=9860 $D=1
M1125 833 137 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=600 $D=1
M1126 834 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=5230 $D=1
M1127 835 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=228150 $Y=9860 $D=1
M1128 836 833 147 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=600 $D=1
M1129 837 834 148 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=5230 $D=1
M1130 838 835 149 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=228885 $Y=9860 $D=1
M1131 141 137 836 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=600 $D=1
M1132 141 137 837 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=5230 $D=1
M1133 141 137 838 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=229405 $Y=9860 $D=1
M1134 839 137 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=600 $D=1
M1135 840 137 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=5230 $D=1
M1136 841 137 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=230140 $Y=9860 $D=1
M1137 842 839 150 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=600 $D=1
M1138 843 840 151 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=5230 $D=1
M1139 844 841 152 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=230875 $Y=9860 $D=1
M1140 141 137 842 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=600 $D=1
M1141 141 137 843 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=5230 $D=1
M1142 141 137 844 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=231395 $Y=9860 $D=1
M1143 7 737 1059 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=600 $D=1
M1144 8 738 1060 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=5230 $D=1
M1145 9 739 1061 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=232130 $Y=9860 $D=1
M1146 142 1059 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=600 $D=1
M1147 138 1060 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=5230 $D=1
M1148 139 1061 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=232510 $Y=9860 $D=1
M1149 845 153 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=600 $D=1
M1150 846 153 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=5230 $D=1
M1151 847 153 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=233170 $Y=9860 $D=1
M1152 146 845 142 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=600 $D=1
M1153 154 846 138 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=5230 $D=1
M1154 143 847 139 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=233905 $Y=9860 $D=1
M1155 818 153 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=600 $D=1
M1156 819 153 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=5230 $D=1
M1157 820 153 143 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=234425 $Y=9860 $D=1
M1158 848 155 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=600 $D=1
M1159 849 155 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=5230 $D=1
M1160 850 155 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=235160 $Y=9860 $D=1
M1161 156 848 146 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=600 $D=1
M1162 157 849 154 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=5230 $D=1
M1163 158 850 143 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=235895 $Y=9860 $D=1
M1164 824 155 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=600 $D=1
M1165 825 155 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=5230 $D=1
M1166 826 155 158 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=236415 $Y=9860 $D=1
M1167 851 159 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=600 $D=1
M1168 852 159 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=5230 $D=1
M1169 853 159 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=237150 $Y=9860 $D=1
M1170 112 851 156 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=600 $D=1
M1171 116 852 157 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=5230 $D=1
M1172 111 853 158 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=237885 $Y=9860 $D=1
M1173 830 159 112 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=600 $D=1
M1174 831 159 116 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=5230 $D=1
M1175 832 159 111 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=238405 $Y=9860 $D=1
M1176 854 160 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=600 $D=1
M1177 855 160 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=5230 $D=1
M1178 856 160 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=239140 $Y=9860 $D=1
M1179 161 854 112 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=600 $D=1
M1180 162 855 116 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=5230 $D=1
M1181 163 856 111 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=239875 $Y=9860 $D=1
M1182 836 160 161 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=600 $D=1
M1183 837 160 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=5230 $D=1
M1184 838 160 163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=240395 $Y=9860 $D=1
M1185 857 164 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=600 $D=1
M1186 858 164 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=5230 $D=1
M1187 859 164 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=241130 $Y=9860 $D=1
M1188 213 857 161 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=600 $D=1
M1189 214 858 162 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=5230 $D=1
M1190 215 859 163 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=241865 $Y=9860 $D=1
M1191 842 164 213 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=600 $D=1
M1192 843 164 214 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=5230 $D=1
M1193 844 164 215 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=242385 $Y=9860 $D=1
M1194 860 165 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=600 $D=1
M1195 861 165 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=5230 $D=1
M1196 862 165 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=243120 $Y=9860 $D=1
M1197 166 860 123 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=600 $D=1
M1198 863 861 124 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=5230 $D=1
M1199 864 862 125 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=243855 $Y=9860 $D=1
M1200 14 165 166 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=600 $D=1
M1201 15 165 863 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=5230 $D=1
M1202 16 165 864 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=244375 $Y=9860 $D=1
M1203 1092 122 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=600 $D=1
M1204 1093 723 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=5230 $D=1
M1205 1094 724 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=9860 $D=1
M1206 865 166 1092 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=600 $D=1
M1207 866 863 1093 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=5230 $D=1
M1208 867 864 1094 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=9860 $D=1
M1209 871 122 868 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=600 $D=1
M1210 872 723 869 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=5230 $D=1
M1211 873 724 870 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=246150 $Y=9860 $D=1
M1212 868 166 871 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=600 $D=1
M1213 869 863 872 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=5230 $D=1
M1214 870 864 873 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.52e-14 PD=6.75e-07 PS=6.4e-07 $X=246530 $Y=9860 $D=1
M1215 7 865 868 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=600 $D=1
M1216 8 866 869 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=5230 $D=1
M1217 9 867 870 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=2.835e-14 PD=6.75e-07 PS=6.75e-07 $X=246945 $Y=9860 $D=1
M1218 1095 167 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=600 $D=1
M1219 1096 874 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=5230 $D=1
M1220 1097 875 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=9860 $D=1
M1221 1062 871 1095 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=600 $D=1
M1222 1063 872 1096 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=5230 $D=1
M1223 1064 873 1097 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=9860 $D=1
M1224 874 1062 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=600 $D=1
M1225 875 1063 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=5230 $D=1
M1226 168 1064 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=248400 $Y=9860 $D=1
M1227 876 122 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=600 $D=1
M1228 877 723 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=5230 $D=1
M1229 878 724 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=249060 $Y=9860 $D=1
M1230 7 879 876 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=600 $D=1
M1231 8 880 877 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=5230 $D=1
M1232 9 881 878 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=249440 $Y=9860 $D=1
M1233 879 166 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=600 $D=1
M1234 880 863 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=5230 $D=1
M1235 881 864 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=250100 $Y=9860 $D=1
M1236 1098 876 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=600 $D=1
M1237 1099 877 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=5230 $D=1
M1238 1100 878 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=9860 $D=1
M1239 882 167 1098 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=600 $D=1
M1240 883 874 1099 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=5230 $D=1
M1241 884 875 1100 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=9860 $D=1
M1242 887 7 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=600 $D=1
M1243 888 885 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=5230 $D=1
M1244 889 886 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=251800 $Y=9860 $D=1
M1245 1101 882 7 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=600 $D=1
M1246 1102 883 8 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=5230 $D=1
M1247 1103 884 9 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=9860 $D=1
M1248 885 887 1101 7 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=600 $D=1
M1249 886 888 1102 8 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=5230 $D=1
M1250 169 889 1103 9 NMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=9860 $D=1
M1251 892 890 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=600 $D=1
M1252 893 891 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=5230 $D=1
M1253 894 170 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=253500 $Y=9860 $D=1
M1254 7 898 895 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=600 $D=1
M1255 8 899 896 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=5230 $D=1
M1256 9 900 897 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=254160 $Y=9860 $D=1
M1257 901 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=600 $D=1
M1258 902 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=5230 $D=1
M1259 903 129 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=254540 $Y=9860 $D=1
M1260 898 901 890 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=600 $D=1
M1261 899 902 891 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=5230 $D=1
M1262 900 903 170 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=255275 $Y=9860 $D=1
M1263 892 127 898 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=600 $D=1
M1264 893 128 899 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=5230 $D=1
M1265 894 129 900 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=255795 $Y=9860 $D=1
M1266 904 895 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=600 $D=1
M1267 905 896 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=5230 $D=1
M1268 906 897 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=256530 $Y=9860 $D=1
M1269 907 904 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=600 $D=1
M1270 890 905 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=5230 $D=1
M1271 891 906 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=257265 $Y=9860 $D=1
M1272 127 895 907 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=600 $D=1
M1273 128 896 890 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=5230 $D=1
M1274 129 897 891 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=257785 $Y=9860 $D=1
M1275 908 907 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=600 $D=1
M1276 909 890 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=5230 $D=1
M1277 910 891 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=258520 $Y=9860 $D=1
M1278 911 895 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=600 $D=1
M1279 912 896 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=5230 $D=1
M1280 913 897 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=259180 $Y=9860 $D=1
M1281 216 911 908 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=600 $D=1
M1282 217 912 909 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=5230 $D=1
M1283 218 913 910 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=259915 $Y=9860 $D=1
M1284 7 895 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=600 $D=1
M1285 8 896 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=5230 $D=1
M1286 9 897 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=260435 $Y=9860 $D=1
M1287 914 171 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=600 $D=1
M1288 915 171 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=5230 $D=1
M1289 916 171 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=261170 $Y=9860 $D=1
M1290 917 914 216 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=600 $D=1
M1291 918 915 217 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=5230 $D=1
M1292 919 916 218 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=261905 $Y=9860 $D=1
M1293 17 171 917 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=600 $D=1
M1294 18 171 918 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=5230 $D=1
M1295 19 171 919 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=262425 $Y=9860 $D=1
M1296 920 172 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=600 $D=1
M1297 921 172 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=5230 $D=1
M1298 922 172 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=263160 $Y=9860 $D=1
M1299 923 920 917 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=600 $D=1
M1300 172 921 918 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=5230 $D=1
M1301 172 922 919 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=263895 $Y=9860 $D=1
M1302 7 172 923 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=600 $D=1
M1303 173 172 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=5230 $D=1
M1304 174 172 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=264415 $Y=9860 $D=1
M1305 924 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=600 $D=1
M1306 925 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=5230 $D=1
M1307 926 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=265150 $Y=9860 $D=1
M1308 7 924 927 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=600 $D=1
M1309 8 925 928 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=5230 $D=1
M1310 9 926 929 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=265810 $Y=9860 $D=1
M1311 930 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=600 $D=1
M1312 931 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=5230 $D=1
M1313 932 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=266190 $Y=9860 $D=1
M1314 933 924 923 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=600 $D=1
M1315 934 925 172 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=5230 $D=1
M1316 935 926 172 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=266925 $Y=9860 $D=1
M1317 7 933 1065 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=600 $D=1
M1318 8 934 1066 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=5230 $D=1
M1319 9 935 1067 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=267660 $Y=9860 $D=1
M1320 936 1065 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=600 $D=1
M1321 937 1066 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=5230 $D=1
M1322 938 1067 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=268040 $Y=9860 $D=1
M1323 933 927 936 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=600 $D=1
M1324 934 928 937 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=5230 $D=1
M1325 935 929 938 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=268485 $Y=9860 $D=1
M1326 939 121 936 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=600 $D=1
M1327 940 121 937 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=5230 $D=1
M1328 941 121 938 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=269295 $Y=9860 $D=1
M1329 7 945 942 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=600 $D=1
M1330 8 946 943 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=5230 $D=1
M1331 9 947 944 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=270030 $Y=9860 $D=1
M1332 945 121 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=600 $D=1
M1333 946 121 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=5230 $D=1
M1334 947 121 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=270410 $Y=9860 $D=1
M1335 1068 939 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=600 $D=1
M1336 1069 940 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=5230 $D=1
M1337 1070 941 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=271070 $Y=9860 $D=1
M1338 948 942 1068 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=600 $D=1
M1339 949 943 1069 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=5230 $D=1
M1340 950 944 1070 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=271515 $Y=9860 $D=1
M1341 7 948 127 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=600 $D=1
M1342 8 949 128 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=5230 $D=1
M1343 9 950 129 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=272250 $Y=9860 $D=1
M1344 1071 127 7 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=600 $D=1
M1345 1072 128 8 8 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=5230 $D=1
M1346 1073 129 9 9 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=272630 $Y=9860 $D=1
M1347 948 945 1071 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=600 $D=1
M1348 949 946 1072 8 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=5230 $D=1
M1349 950 947 1073 9 NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=273010 $Y=9860 $D=1
M1350 177 1 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M1351 178 1 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=6480 $D=0
M1352 179 1 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=11110 $D=0
M1353 180 1 2 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=1850 $D=0
M1354 181 1 3 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=6480 $D=0
M1355 182 1 4 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=1045 $Y=11110 $D=0
M1356 7 177 180 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=1850 $D=0
M1357 8 178 181 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=6480 $D=0
M1358 9 179 182 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=1565 $Y=11110 $D=0
M1359 183 1 5 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=1850 $D=0
M1360 184 1 5 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=6480 $D=0
M1361 185 1 5 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=2375 $Y=11110 $D=0
M1362 6 177 183 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=1850 $D=0
M1363 6 178 184 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=6480 $D=0
M1364 6 179 185 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=2895 $Y=11110 $D=0
M1365 186 1 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=1850 $D=0
M1366 187 1 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=6480 $D=0
M1367 188 1 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3705 $Y=11110 $D=0
M1368 7 177 186 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=1850 $D=0
M1369 8 178 187 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=6480 $D=0
M1370 9 179 188 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4225 $Y=11110 $D=0
M1371 192 11 186 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=1850 $D=0
M1372 193 11 187 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=6480 $D=0
M1373 194 11 188 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=5035 $Y=11110 $D=0
M1374 189 11 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=1850 $D=0
M1375 190 11 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=6480 $D=0
M1376 191 11 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5770 $Y=11110 $D=0
M1377 195 11 183 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=1850 $D=0
M1378 196 11 184 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=6480 $D=0
M1379 197 11 185 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=6505 $Y=11110 $D=0
M1380 180 189 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=1850 $D=0
M1381 181 190 196 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=6480 $D=0
M1382 182 191 197 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=7025 $Y=11110 $D=0
M1383 198 12 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=1850 $D=0
M1384 199 12 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=6480 $D=0
M1385 200 12 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=7760 $Y=11110 $D=0
M1386 201 12 195 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=1850 $D=0
M1387 202 12 196 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=6480 $D=0
M1388 203 12 197 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=8495 $Y=11110 $D=0
M1389 192 198 201 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=1850 $D=0
M1390 193 199 202 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=6480 $D=0
M1391 194 200 203 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=9015 $Y=11110 $D=0
M1392 204 13 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=1850 $D=0
M1393 205 13 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=6480 $D=0
M1394 206 13 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=9750 $Y=11110 $D=0
M1395 207 13 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=1850 $D=0
M1396 208 13 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=6480 $D=0
M1397 209 13 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=10485 $Y=11110 $D=0
M1398 14 204 207 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=1850 $D=0
M1399 15 205 208 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=6480 $D=0
M1400 16 206 209 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=11005 $Y=11110 $D=0
M1401 210 13 17 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=1850 $D=0
M1402 211 13 18 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=6480 $D=0
M1403 212 13 19 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=11815 $Y=11110 $D=0
M1404 213 204 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=1850 $D=0
M1405 214 205 211 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=6480 $D=0
M1406 215 206 212 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=12335 $Y=11110 $D=0
M1407 219 13 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=1850 $D=0
M1408 220 13 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=6480 $D=0
M1409 221 13 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=13145 $Y=11110 $D=0
M1410 201 204 219 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=1850 $D=0
M1411 202 205 220 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=6480 $D=0
M1412 203 206 221 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=13665 $Y=11110 $D=0
M1413 225 20 219 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=1850 $D=0
M1414 226 20 220 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=6480 $D=0
M1415 227 20 221 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=14475 $Y=11110 $D=0
M1416 222 20 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=1850 $D=0
M1417 223 20 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=6480 $D=0
M1418 224 20 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=15210 $Y=11110 $D=0
M1419 228 20 210 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=1850 $D=0
M1420 229 20 211 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=6480 $D=0
M1421 230 20 212 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=15945 $Y=11110 $D=0
M1422 207 222 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=1850 $D=0
M1423 208 223 229 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=6480 $D=0
M1424 209 224 230 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=16465 $Y=11110 $D=0
M1425 231 21 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=1850 $D=0
M1426 232 21 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=6480 $D=0
M1427 233 21 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=17200 $Y=11110 $D=0
M1428 234 21 228 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=1850 $D=0
M1429 235 21 229 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=6480 $D=0
M1430 236 21 230 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=17935 $Y=11110 $D=0
M1431 225 231 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=1850 $D=0
M1432 226 232 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=6480 $D=0
M1433 227 233 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=18455 $Y=11110 $D=0
M1434 167 22 237 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=1850 $D=0
M1435 173 22 238 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=6480 $D=0
M1436 174 22 239 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=19190 $Y=11110 $D=0
M1437 240 23 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=1850 $D=0
M1438 241 23 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=6480 $D=0
M1439 242 23 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=19570 $Y=11110 $D=0
M1440 243 237 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=1850 $D=0
M1441 244 238 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=6480 $D=0
M1442 245 239 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=20305 $Y=11110 $D=0
M1443 167 243 951 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=1850 $D=0
M1444 173 244 952 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=6480 $D=0
M1445 174 245 953 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=21040 $Y=11110 $D=0
M1446 246 951 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=1850 $D=0
M1447 247 952 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=6480 $D=0
M1448 248 953 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=21420 $Y=11110 $D=0
M1449 243 22 246 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=1850 $D=0
M1450 244 22 247 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=6480 $D=0
M1451 245 22 248 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=21865 $Y=11110 $D=0
M1452 246 240 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=1850 $D=0
M1453 247 241 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=6480 $D=0
M1454 248 242 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=22675 $Y=11110 $D=0
M1455 255 252 246 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=1850 $D=0
M1456 256 253 247 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=6480 $D=0
M1457 257 254 248 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=23195 $Y=11110 $D=0
M1458 252 24 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=1850 $D=0
M1459 253 24 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=6480 $D=0
M1460 254 24 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=23930 $Y=11110 $D=0
M1461 167 25 258 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=1850 $D=0
M1462 173 25 259 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=6480 $D=0
M1463 174 25 260 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=24590 $Y=11110 $D=0
M1464 261 26 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=1850 $D=0
M1465 262 26 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=6480 $D=0
M1466 263 26 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=24970 $Y=11110 $D=0
M1467 264 258 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=1850 $D=0
M1468 265 259 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=6480 $D=0
M1469 266 260 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=25705 $Y=11110 $D=0
M1470 167 264 954 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=1850 $D=0
M1471 173 265 955 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=6480 $D=0
M1472 174 266 956 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=26440 $Y=11110 $D=0
M1473 267 954 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=1850 $D=0
M1474 268 955 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=6480 $D=0
M1475 269 956 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=26820 $Y=11110 $D=0
M1476 264 25 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=1850 $D=0
M1477 265 25 268 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=6480 $D=0
M1478 266 25 269 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=27265 $Y=11110 $D=0
M1479 267 261 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=1850 $D=0
M1480 268 262 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=6480 $D=0
M1481 269 263 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=28075 $Y=11110 $D=0
M1482 255 270 267 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=1850 $D=0
M1483 256 271 268 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=6480 $D=0
M1484 257 272 269 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=28595 $Y=11110 $D=0
M1485 270 27 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=1850 $D=0
M1486 271 27 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=6480 $D=0
M1487 272 27 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=29330 $Y=11110 $D=0
M1488 167 28 273 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=1850 $D=0
M1489 173 28 274 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=6480 $D=0
M1490 174 28 275 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=29990 $Y=11110 $D=0
M1491 276 29 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=1850 $D=0
M1492 277 29 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=6480 $D=0
M1493 278 29 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=30370 $Y=11110 $D=0
M1494 279 273 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=1850 $D=0
M1495 280 274 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=6480 $D=0
M1496 281 275 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=31105 $Y=11110 $D=0
M1497 167 279 957 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=1850 $D=0
M1498 173 280 958 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=6480 $D=0
M1499 174 281 959 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=31840 $Y=11110 $D=0
M1500 282 957 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=1850 $D=0
M1501 283 958 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=6480 $D=0
M1502 284 959 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=32220 $Y=11110 $D=0
M1503 279 28 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=1850 $D=0
M1504 280 28 283 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=6480 $D=0
M1505 281 28 284 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=32665 $Y=11110 $D=0
M1506 282 276 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=1850 $D=0
M1507 283 277 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=6480 $D=0
M1508 284 278 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=33475 $Y=11110 $D=0
M1509 255 285 282 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=1850 $D=0
M1510 256 286 283 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=6480 $D=0
M1511 257 287 284 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=33995 $Y=11110 $D=0
M1512 285 30 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=1850 $D=0
M1513 286 30 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=6480 $D=0
M1514 287 30 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=34730 $Y=11110 $D=0
M1515 167 31 288 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=1850 $D=0
M1516 173 31 289 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=6480 $D=0
M1517 174 31 290 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=35390 $Y=11110 $D=0
M1518 291 32 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=1850 $D=0
M1519 292 32 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=6480 $D=0
M1520 293 32 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=35770 $Y=11110 $D=0
M1521 294 288 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=1850 $D=0
M1522 295 289 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=6480 $D=0
M1523 296 290 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=36505 $Y=11110 $D=0
M1524 167 294 960 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=1850 $D=0
M1525 173 295 961 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=6480 $D=0
M1526 174 296 962 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=37240 $Y=11110 $D=0
M1527 297 960 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=1850 $D=0
M1528 298 961 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=6480 $D=0
M1529 299 962 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=37620 $Y=11110 $D=0
M1530 294 31 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=1850 $D=0
M1531 295 31 298 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=6480 $D=0
M1532 296 31 299 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=38065 $Y=11110 $D=0
M1533 297 291 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=1850 $D=0
M1534 298 292 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=6480 $D=0
M1535 299 293 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=38875 $Y=11110 $D=0
M1536 255 300 297 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=1850 $D=0
M1537 256 301 298 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=6480 $D=0
M1538 257 302 299 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=39395 $Y=11110 $D=0
M1539 300 33 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=1850 $D=0
M1540 301 33 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=6480 $D=0
M1541 302 33 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=40130 $Y=11110 $D=0
M1542 167 34 303 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=1850 $D=0
M1543 173 34 304 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=6480 $D=0
M1544 174 34 305 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=40790 $Y=11110 $D=0
M1545 306 35 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=1850 $D=0
M1546 307 35 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=6480 $D=0
M1547 308 35 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=41170 $Y=11110 $D=0
M1548 309 303 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=1850 $D=0
M1549 310 304 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=6480 $D=0
M1550 311 305 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=41905 $Y=11110 $D=0
M1551 167 309 963 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=1850 $D=0
M1552 173 310 964 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=6480 $D=0
M1553 174 311 965 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=42640 $Y=11110 $D=0
M1554 312 963 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=1850 $D=0
M1555 313 964 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=6480 $D=0
M1556 314 965 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=43020 $Y=11110 $D=0
M1557 309 34 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=1850 $D=0
M1558 310 34 313 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=6480 $D=0
M1559 311 34 314 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=43465 $Y=11110 $D=0
M1560 312 306 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=1850 $D=0
M1561 313 307 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=6480 $D=0
M1562 314 308 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=44275 $Y=11110 $D=0
M1563 255 315 312 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=1850 $D=0
M1564 256 316 313 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=6480 $D=0
M1565 257 317 314 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=44795 $Y=11110 $D=0
M1566 315 36 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=1850 $D=0
M1567 316 36 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=6480 $D=0
M1568 317 36 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=45530 $Y=11110 $D=0
M1569 167 37 318 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=1850 $D=0
M1570 173 37 319 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=6480 $D=0
M1571 174 37 320 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=46190 $Y=11110 $D=0
M1572 321 38 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=1850 $D=0
M1573 322 38 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=6480 $D=0
M1574 323 38 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=46570 $Y=11110 $D=0
M1575 324 318 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=1850 $D=0
M1576 325 319 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=6480 $D=0
M1577 326 320 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=47305 $Y=11110 $D=0
M1578 167 324 966 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=1850 $D=0
M1579 173 325 967 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=6480 $D=0
M1580 174 326 968 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=48040 $Y=11110 $D=0
M1581 327 966 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=1850 $D=0
M1582 328 967 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=6480 $D=0
M1583 329 968 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=48420 $Y=11110 $D=0
M1584 324 37 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=1850 $D=0
M1585 325 37 328 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=6480 $D=0
M1586 326 37 329 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=48865 $Y=11110 $D=0
M1587 327 321 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=1850 $D=0
M1588 328 322 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=6480 $D=0
M1589 329 323 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=49675 $Y=11110 $D=0
M1590 255 330 327 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=1850 $D=0
M1591 256 331 328 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=6480 $D=0
M1592 257 332 329 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=50195 $Y=11110 $D=0
M1593 330 39 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=1850 $D=0
M1594 331 39 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=6480 $D=0
M1595 332 39 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=50930 $Y=11110 $D=0
M1596 167 40 333 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=1850 $D=0
M1597 173 40 334 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=6480 $D=0
M1598 174 40 335 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=51590 $Y=11110 $D=0
M1599 336 41 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=1850 $D=0
M1600 337 41 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=6480 $D=0
M1601 338 41 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=51970 $Y=11110 $D=0
M1602 339 333 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=1850 $D=0
M1603 340 334 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=6480 $D=0
M1604 341 335 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=52705 $Y=11110 $D=0
M1605 167 339 969 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=1850 $D=0
M1606 173 340 970 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=6480 $D=0
M1607 174 341 971 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=53440 $Y=11110 $D=0
M1608 342 969 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=1850 $D=0
M1609 343 970 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=6480 $D=0
M1610 344 971 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=53820 $Y=11110 $D=0
M1611 339 40 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=1850 $D=0
M1612 340 40 343 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=6480 $D=0
M1613 341 40 344 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=54265 $Y=11110 $D=0
M1614 342 336 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=1850 $D=0
M1615 343 337 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=6480 $D=0
M1616 344 338 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=55075 $Y=11110 $D=0
M1617 255 345 342 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=1850 $D=0
M1618 256 346 343 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=6480 $D=0
M1619 257 347 344 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=55595 $Y=11110 $D=0
M1620 345 42 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=1850 $D=0
M1621 346 42 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=6480 $D=0
M1622 347 42 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=56330 $Y=11110 $D=0
M1623 167 43 348 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=1850 $D=0
M1624 173 43 349 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=6480 $D=0
M1625 174 43 350 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=56990 $Y=11110 $D=0
M1626 351 44 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=1850 $D=0
M1627 352 44 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=6480 $D=0
M1628 353 44 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=57370 $Y=11110 $D=0
M1629 354 348 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=1850 $D=0
M1630 355 349 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=6480 $D=0
M1631 356 350 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=58105 $Y=11110 $D=0
M1632 167 354 972 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=1850 $D=0
M1633 173 355 973 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=6480 $D=0
M1634 174 356 974 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=58840 $Y=11110 $D=0
M1635 357 972 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=1850 $D=0
M1636 358 973 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=6480 $D=0
M1637 359 974 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=59220 $Y=11110 $D=0
M1638 354 43 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=1850 $D=0
M1639 355 43 358 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=6480 $D=0
M1640 356 43 359 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=59665 $Y=11110 $D=0
M1641 357 351 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=1850 $D=0
M1642 358 352 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=6480 $D=0
M1643 359 353 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=60475 $Y=11110 $D=0
M1644 255 360 357 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=1850 $D=0
M1645 256 361 358 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=6480 $D=0
M1646 257 362 359 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=60995 $Y=11110 $D=0
M1647 360 45 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=1850 $D=0
M1648 361 45 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=6480 $D=0
M1649 362 45 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=61730 $Y=11110 $D=0
M1650 167 46 363 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=1850 $D=0
M1651 173 46 364 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=6480 $D=0
M1652 174 46 365 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=62390 $Y=11110 $D=0
M1653 366 47 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=1850 $D=0
M1654 367 47 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=6480 $D=0
M1655 368 47 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=62770 $Y=11110 $D=0
M1656 369 363 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=1850 $D=0
M1657 370 364 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=6480 $D=0
M1658 371 365 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=63505 $Y=11110 $D=0
M1659 167 369 975 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=1850 $D=0
M1660 173 370 976 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=6480 $D=0
M1661 174 371 977 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=64240 $Y=11110 $D=0
M1662 372 975 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=1850 $D=0
M1663 373 976 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=6480 $D=0
M1664 374 977 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=64620 $Y=11110 $D=0
M1665 369 46 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=1850 $D=0
M1666 370 46 373 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=6480 $D=0
M1667 371 46 374 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=65065 $Y=11110 $D=0
M1668 372 366 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=1850 $D=0
M1669 373 367 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=6480 $D=0
M1670 374 368 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=65875 $Y=11110 $D=0
M1671 255 375 372 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=1850 $D=0
M1672 256 376 373 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=6480 $D=0
M1673 257 377 374 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=66395 $Y=11110 $D=0
M1674 375 48 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=1850 $D=0
M1675 376 48 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=6480 $D=0
M1676 377 48 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=67130 $Y=11110 $D=0
M1677 167 49 378 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=1850 $D=0
M1678 173 49 379 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=6480 $D=0
M1679 174 49 380 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=67790 $Y=11110 $D=0
M1680 381 50 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=1850 $D=0
M1681 382 50 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=6480 $D=0
M1682 383 50 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=68170 $Y=11110 $D=0
M1683 384 378 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=1850 $D=0
M1684 385 379 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=6480 $D=0
M1685 386 380 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=68905 $Y=11110 $D=0
M1686 167 384 978 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=1850 $D=0
M1687 173 385 979 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=6480 $D=0
M1688 174 386 980 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=69640 $Y=11110 $D=0
M1689 387 978 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=1850 $D=0
M1690 388 979 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=6480 $D=0
M1691 389 980 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=70020 $Y=11110 $D=0
M1692 384 49 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=1850 $D=0
M1693 385 49 388 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=6480 $D=0
M1694 386 49 389 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=70465 $Y=11110 $D=0
M1695 387 381 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=1850 $D=0
M1696 388 382 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=6480 $D=0
M1697 389 383 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=71275 $Y=11110 $D=0
M1698 255 390 387 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=1850 $D=0
M1699 256 391 388 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=6480 $D=0
M1700 257 392 389 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=71795 $Y=11110 $D=0
M1701 390 51 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=1850 $D=0
M1702 391 51 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=6480 $D=0
M1703 392 51 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=72530 $Y=11110 $D=0
M1704 167 52 393 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=1850 $D=0
M1705 173 52 394 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=6480 $D=0
M1706 174 52 395 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=73190 $Y=11110 $D=0
M1707 396 53 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=1850 $D=0
M1708 397 53 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=6480 $D=0
M1709 398 53 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=73570 $Y=11110 $D=0
M1710 399 393 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=1850 $D=0
M1711 400 394 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=6480 $D=0
M1712 401 395 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=74305 $Y=11110 $D=0
M1713 167 399 981 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=1850 $D=0
M1714 173 400 982 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=6480 $D=0
M1715 174 401 983 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=75040 $Y=11110 $D=0
M1716 402 981 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=1850 $D=0
M1717 403 982 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=6480 $D=0
M1718 404 983 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=75420 $Y=11110 $D=0
M1719 399 52 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=1850 $D=0
M1720 400 52 403 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=6480 $D=0
M1721 401 52 404 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=75865 $Y=11110 $D=0
M1722 402 396 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=1850 $D=0
M1723 403 397 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=6480 $D=0
M1724 404 398 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=76675 $Y=11110 $D=0
M1725 255 405 402 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=1850 $D=0
M1726 256 406 403 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=6480 $D=0
M1727 257 407 404 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=77195 $Y=11110 $D=0
M1728 405 54 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=1850 $D=0
M1729 406 54 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=6480 $D=0
M1730 407 54 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=77930 $Y=11110 $D=0
M1731 167 55 408 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=1850 $D=0
M1732 173 55 409 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=6480 $D=0
M1733 174 55 410 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=78590 $Y=11110 $D=0
M1734 411 56 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=1850 $D=0
M1735 412 56 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=6480 $D=0
M1736 413 56 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=78970 $Y=11110 $D=0
M1737 414 408 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=1850 $D=0
M1738 415 409 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=6480 $D=0
M1739 416 410 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=79705 $Y=11110 $D=0
M1740 167 414 984 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=1850 $D=0
M1741 173 415 985 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=6480 $D=0
M1742 174 416 986 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=80440 $Y=11110 $D=0
M1743 417 984 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=1850 $D=0
M1744 418 985 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=6480 $D=0
M1745 419 986 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=80820 $Y=11110 $D=0
M1746 414 55 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=1850 $D=0
M1747 415 55 418 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=6480 $D=0
M1748 416 55 419 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=81265 $Y=11110 $D=0
M1749 417 411 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=1850 $D=0
M1750 418 412 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=6480 $D=0
M1751 419 413 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=82075 $Y=11110 $D=0
M1752 255 420 417 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=1850 $D=0
M1753 256 421 418 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=6480 $D=0
M1754 257 422 419 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=82595 $Y=11110 $D=0
M1755 420 57 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=1850 $D=0
M1756 421 57 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=6480 $D=0
M1757 422 57 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=83330 $Y=11110 $D=0
M1758 167 58 423 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=1850 $D=0
M1759 173 58 424 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=6480 $D=0
M1760 174 58 425 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=83990 $Y=11110 $D=0
M1761 426 59 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=1850 $D=0
M1762 427 59 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=6480 $D=0
M1763 428 59 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=84370 $Y=11110 $D=0
M1764 429 423 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=1850 $D=0
M1765 430 424 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=6480 $D=0
M1766 431 425 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=85105 $Y=11110 $D=0
M1767 167 429 987 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=1850 $D=0
M1768 173 430 988 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=6480 $D=0
M1769 174 431 989 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=85840 $Y=11110 $D=0
M1770 432 987 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=1850 $D=0
M1771 433 988 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=6480 $D=0
M1772 434 989 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=86220 $Y=11110 $D=0
M1773 429 58 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=1850 $D=0
M1774 430 58 433 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=6480 $D=0
M1775 431 58 434 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=86665 $Y=11110 $D=0
M1776 432 426 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=1850 $D=0
M1777 433 427 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=6480 $D=0
M1778 434 428 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=87475 $Y=11110 $D=0
M1779 255 435 432 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=1850 $D=0
M1780 256 436 433 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=6480 $D=0
M1781 257 437 434 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=87995 $Y=11110 $D=0
M1782 435 60 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=1850 $D=0
M1783 436 60 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=6480 $D=0
M1784 437 60 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=88730 $Y=11110 $D=0
M1785 167 61 438 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=1850 $D=0
M1786 173 61 439 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=6480 $D=0
M1787 174 61 440 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=89390 $Y=11110 $D=0
M1788 441 62 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=1850 $D=0
M1789 442 62 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=6480 $D=0
M1790 443 62 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=89770 $Y=11110 $D=0
M1791 444 438 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=1850 $D=0
M1792 445 439 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=6480 $D=0
M1793 446 440 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=90505 $Y=11110 $D=0
M1794 167 444 990 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=1850 $D=0
M1795 173 445 991 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=6480 $D=0
M1796 174 446 992 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=91240 $Y=11110 $D=0
M1797 447 990 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=1850 $D=0
M1798 448 991 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=6480 $D=0
M1799 449 992 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=91620 $Y=11110 $D=0
M1800 444 61 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=1850 $D=0
M1801 445 61 448 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=6480 $D=0
M1802 446 61 449 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=92065 $Y=11110 $D=0
M1803 447 441 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=1850 $D=0
M1804 448 442 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=6480 $D=0
M1805 449 443 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=92875 $Y=11110 $D=0
M1806 255 450 447 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=1850 $D=0
M1807 256 451 448 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=6480 $D=0
M1808 257 452 449 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=93395 $Y=11110 $D=0
M1809 450 63 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=1850 $D=0
M1810 451 63 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=6480 $D=0
M1811 452 63 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=94130 $Y=11110 $D=0
M1812 167 64 453 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=1850 $D=0
M1813 173 64 454 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=6480 $D=0
M1814 174 64 455 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=94790 $Y=11110 $D=0
M1815 456 65 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=1850 $D=0
M1816 457 65 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=6480 $D=0
M1817 458 65 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=95170 $Y=11110 $D=0
M1818 459 453 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=1850 $D=0
M1819 460 454 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=6480 $D=0
M1820 461 455 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=95905 $Y=11110 $D=0
M1821 167 459 993 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=1850 $D=0
M1822 173 460 994 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=6480 $D=0
M1823 174 461 995 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=96640 $Y=11110 $D=0
M1824 462 993 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=1850 $D=0
M1825 463 994 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=6480 $D=0
M1826 464 995 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=97020 $Y=11110 $D=0
M1827 459 64 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=1850 $D=0
M1828 460 64 463 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=6480 $D=0
M1829 461 64 464 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=97465 $Y=11110 $D=0
M1830 462 456 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=1850 $D=0
M1831 463 457 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=6480 $D=0
M1832 464 458 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=98275 $Y=11110 $D=0
M1833 255 465 462 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=1850 $D=0
M1834 256 466 463 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=6480 $D=0
M1835 257 467 464 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=98795 $Y=11110 $D=0
M1836 465 66 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=1850 $D=0
M1837 466 66 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=6480 $D=0
M1838 467 66 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=99530 $Y=11110 $D=0
M1839 167 67 468 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=1850 $D=0
M1840 173 67 469 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=6480 $D=0
M1841 174 67 470 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=100190 $Y=11110 $D=0
M1842 471 68 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=1850 $D=0
M1843 472 68 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=6480 $D=0
M1844 473 68 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=100570 $Y=11110 $D=0
M1845 474 468 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=1850 $D=0
M1846 475 469 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=6480 $D=0
M1847 476 470 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=101305 $Y=11110 $D=0
M1848 167 474 996 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=1850 $D=0
M1849 173 475 997 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=6480 $D=0
M1850 174 476 998 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=102040 $Y=11110 $D=0
M1851 477 996 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=1850 $D=0
M1852 478 997 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=6480 $D=0
M1853 479 998 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=102420 $Y=11110 $D=0
M1854 474 67 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=1850 $D=0
M1855 475 67 478 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=6480 $D=0
M1856 476 67 479 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=102865 $Y=11110 $D=0
M1857 477 471 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=1850 $D=0
M1858 478 472 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=6480 $D=0
M1859 479 473 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=103675 $Y=11110 $D=0
M1860 255 480 477 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=1850 $D=0
M1861 256 481 478 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=6480 $D=0
M1862 257 482 479 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=104195 $Y=11110 $D=0
M1863 480 69 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=1850 $D=0
M1864 481 69 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=6480 $D=0
M1865 482 69 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=104930 $Y=11110 $D=0
M1866 167 70 483 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=1850 $D=0
M1867 173 70 484 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=6480 $D=0
M1868 174 70 485 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=105590 $Y=11110 $D=0
M1869 486 71 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=1850 $D=0
M1870 487 71 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=6480 $D=0
M1871 488 71 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=105970 $Y=11110 $D=0
M1872 489 483 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=1850 $D=0
M1873 490 484 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=6480 $D=0
M1874 491 485 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=106705 $Y=11110 $D=0
M1875 167 489 999 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=1850 $D=0
M1876 173 490 1000 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=6480 $D=0
M1877 174 491 1001 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=107440 $Y=11110 $D=0
M1878 492 999 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=1850 $D=0
M1879 493 1000 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=6480 $D=0
M1880 494 1001 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=107820 $Y=11110 $D=0
M1881 489 70 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=1850 $D=0
M1882 490 70 493 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=6480 $D=0
M1883 491 70 494 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=108265 $Y=11110 $D=0
M1884 492 486 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=1850 $D=0
M1885 493 487 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=6480 $D=0
M1886 494 488 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=109075 $Y=11110 $D=0
M1887 255 495 492 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=1850 $D=0
M1888 256 496 493 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=6480 $D=0
M1889 257 497 494 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=109595 $Y=11110 $D=0
M1890 495 72 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=1850 $D=0
M1891 496 72 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=6480 $D=0
M1892 497 72 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=110330 $Y=11110 $D=0
M1893 167 73 498 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=1850 $D=0
M1894 173 73 499 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=6480 $D=0
M1895 174 73 500 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=110990 $Y=11110 $D=0
M1896 501 74 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=1850 $D=0
M1897 502 74 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=6480 $D=0
M1898 503 74 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=111370 $Y=11110 $D=0
M1899 504 498 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=1850 $D=0
M1900 505 499 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=6480 $D=0
M1901 506 500 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=112105 $Y=11110 $D=0
M1902 167 504 1002 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=1850 $D=0
M1903 173 505 1003 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=6480 $D=0
M1904 174 506 1004 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=112840 $Y=11110 $D=0
M1905 507 1002 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=1850 $D=0
M1906 508 1003 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=6480 $D=0
M1907 509 1004 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=113220 $Y=11110 $D=0
M1908 504 73 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=1850 $D=0
M1909 505 73 508 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=6480 $D=0
M1910 506 73 509 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=113665 $Y=11110 $D=0
M1911 507 501 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=1850 $D=0
M1912 508 502 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=6480 $D=0
M1913 509 503 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=114475 $Y=11110 $D=0
M1914 255 510 507 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=1850 $D=0
M1915 256 511 508 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=6480 $D=0
M1916 257 512 509 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=114995 $Y=11110 $D=0
M1917 510 75 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=1850 $D=0
M1918 511 75 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=6480 $D=0
M1919 512 75 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=115730 $Y=11110 $D=0
M1920 167 76 513 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=1850 $D=0
M1921 173 76 514 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=6480 $D=0
M1922 174 76 515 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=116390 $Y=11110 $D=0
M1923 516 77 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=1850 $D=0
M1924 517 77 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=6480 $D=0
M1925 518 77 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=116770 $Y=11110 $D=0
M1926 519 513 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=1850 $D=0
M1927 520 514 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=6480 $D=0
M1928 521 515 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=117505 $Y=11110 $D=0
M1929 167 519 1005 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=1850 $D=0
M1930 173 520 1006 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=6480 $D=0
M1931 174 521 1007 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=118240 $Y=11110 $D=0
M1932 522 1005 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=1850 $D=0
M1933 523 1006 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=6480 $D=0
M1934 524 1007 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=118620 $Y=11110 $D=0
M1935 519 76 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=1850 $D=0
M1936 520 76 523 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=6480 $D=0
M1937 521 76 524 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=119065 $Y=11110 $D=0
M1938 522 516 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=1850 $D=0
M1939 523 517 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=6480 $D=0
M1940 524 518 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=119875 $Y=11110 $D=0
M1941 255 525 522 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=1850 $D=0
M1942 256 526 523 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=6480 $D=0
M1943 257 527 524 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=120395 $Y=11110 $D=0
M1944 525 78 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=1850 $D=0
M1945 526 78 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=6480 $D=0
M1946 527 78 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=121130 $Y=11110 $D=0
M1947 167 79 528 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=1850 $D=0
M1948 173 79 529 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=6480 $D=0
M1949 174 79 530 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=121790 $Y=11110 $D=0
M1950 531 80 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=1850 $D=0
M1951 532 80 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=6480 $D=0
M1952 533 80 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=122170 $Y=11110 $D=0
M1953 534 528 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=1850 $D=0
M1954 535 529 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=6480 $D=0
M1955 536 530 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=122905 $Y=11110 $D=0
M1956 167 534 1008 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=1850 $D=0
M1957 173 535 1009 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=6480 $D=0
M1958 174 536 1010 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=123640 $Y=11110 $D=0
M1959 537 1008 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=1850 $D=0
M1960 538 1009 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=6480 $D=0
M1961 539 1010 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=124020 $Y=11110 $D=0
M1962 534 79 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=1850 $D=0
M1963 535 79 538 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=6480 $D=0
M1964 536 79 539 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=124465 $Y=11110 $D=0
M1965 537 531 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=1850 $D=0
M1966 538 532 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=6480 $D=0
M1967 539 533 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=125275 $Y=11110 $D=0
M1968 255 540 537 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=1850 $D=0
M1969 256 541 538 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=6480 $D=0
M1970 257 542 539 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=125795 $Y=11110 $D=0
M1971 540 81 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=1850 $D=0
M1972 541 81 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=6480 $D=0
M1973 542 81 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=126530 $Y=11110 $D=0
M1974 167 82 543 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=1850 $D=0
M1975 173 82 544 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=6480 $D=0
M1976 174 82 545 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=127190 $Y=11110 $D=0
M1977 546 83 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=1850 $D=0
M1978 547 83 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=6480 $D=0
M1979 548 83 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=127570 $Y=11110 $D=0
M1980 549 543 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=1850 $D=0
M1981 550 544 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=6480 $D=0
M1982 551 545 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=128305 $Y=11110 $D=0
M1983 167 549 1011 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=1850 $D=0
M1984 173 550 1012 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=6480 $D=0
M1985 174 551 1013 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=129040 $Y=11110 $D=0
M1986 552 1011 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=1850 $D=0
M1987 553 1012 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=6480 $D=0
M1988 554 1013 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=129420 $Y=11110 $D=0
M1989 549 82 552 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=1850 $D=0
M1990 550 82 553 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=6480 $D=0
M1991 551 82 554 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=129865 $Y=11110 $D=0
M1992 552 546 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=1850 $D=0
M1993 553 547 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=6480 $D=0
M1994 554 548 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=130675 $Y=11110 $D=0
M1995 255 555 552 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=1850 $D=0
M1996 256 556 553 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=6480 $D=0
M1997 257 557 554 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=131195 $Y=11110 $D=0
M1998 555 84 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=1850 $D=0
M1999 556 84 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=6480 $D=0
M2000 557 84 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=131930 $Y=11110 $D=0
M2001 167 85 558 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=1850 $D=0
M2002 173 85 559 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=6480 $D=0
M2003 174 85 560 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=132590 $Y=11110 $D=0
M2004 561 86 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=1850 $D=0
M2005 562 86 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=6480 $D=0
M2006 563 86 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=132970 $Y=11110 $D=0
M2007 564 558 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=1850 $D=0
M2008 565 559 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=6480 $D=0
M2009 566 560 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=133705 $Y=11110 $D=0
M2010 167 564 1014 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=1850 $D=0
M2011 173 565 1015 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=6480 $D=0
M2012 174 566 1016 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=134440 $Y=11110 $D=0
M2013 567 1014 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=1850 $D=0
M2014 568 1015 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=6480 $D=0
M2015 569 1016 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=134820 $Y=11110 $D=0
M2016 564 85 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=1850 $D=0
M2017 565 85 568 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=6480 $D=0
M2018 566 85 569 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=135265 $Y=11110 $D=0
M2019 567 561 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=1850 $D=0
M2020 568 562 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=6480 $D=0
M2021 569 563 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=136075 $Y=11110 $D=0
M2022 255 570 567 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=1850 $D=0
M2023 256 571 568 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=6480 $D=0
M2024 257 572 569 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=136595 $Y=11110 $D=0
M2025 570 87 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=1850 $D=0
M2026 571 87 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=6480 $D=0
M2027 572 87 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=137330 $Y=11110 $D=0
M2028 167 88 573 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=1850 $D=0
M2029 173 88 574 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=6480 $D=0
M2030 174 88 575 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=137990 $Y=11110 $D=0
M2031 576 89 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=1850 $D=0
M2032 577 89 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=6480 $D=0
M2033 578 89 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=138370 $Y=11110 $D=0
M2034 579 573 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=1850 $D=0
M2035 580 574 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=6480 $D=0
M2036 581 575 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=139105 $Y=11110 $D=0
M2037 167 579 1017 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=1850 $D=0
M2038 173 580 1018 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=6480 $D=0
M2039 174 581 1019 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=139840 $Y=11110 $D=0
M2040 582 1017 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=1850 $D=0
M2041 583 1018 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=6480 $D=0
M2042 584 1019 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=140220 $Y=11110 $D=0
M2043 579 88 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=1850 $D=0
M2044 580 88 583 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=6480 $D=0
M2045 581 88 584 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=140665 $Y=11110 $D=0
M2046 582 576 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=1850 $D=0
M2047 583 577 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=6480 $D=0
M2048 584 578 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=141475 $Y=11110 $D=0
M2049 255 585 582 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=1850 $D=0
M2050 256 586 583 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=6480 $D=0
M2051 257 587 584 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=141995 $Y=11110 $D=0
M2052 585 90 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=1850 $D=0
M2053 586 90 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=6480 $D=0
M2054 587 90 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=142730 $Y=11110 $D=0
M2055 167 91 588 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=1850 $D=0
M2056 173 91 589 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=6480 $D=0
M2057 174 91 590 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=143390 $Y=11110 $D=0
M2058 591 92 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=1850 $D=0
M2059 592 92 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=6480 $D=0
M2060 593 92 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=143770 $Y=11110 $D=0
M2061 594 588 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=1850 $D=0
M2062 595 589 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=6480 $D=0
M2063 596 590 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=144505 $Y=11110 $D=0
M2064 167 594 1020 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=1850 $D=0
M2065 173 595 1021 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=6480 $D=0
M2066 174 596 1022 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=145240 $Y=11110 $D=0
M2067 597 1020 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=1850 $D=0
M2068 598 1021 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=6480 $D=0
M2069 599 1022 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=145620 $Y=11110 $D=0
M2070 594 91 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=1850 $D=0
M2071 595 91 598 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=6480 $D=0
M2072 596 91 599 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=146065 $Y=11110 $D=0
M2073 597 591 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=1850 $D=0
M2074 598 592 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=6480 $D=0
M2075 599 593 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=146875 $Y=11110 $D=0
M2076 255 600 597 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=1850 $D=0
M2077 256 601 598 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=6480 $D=0
M2078 257 602 599 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=147395 $Y=11110 $D=0
M2079 600 93 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=1850 $D=0
M2080 601 93 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=6480 $D=0
M2081 602 93 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=148130 $Y=11110 $D=0
M2082 167 94 603 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=1850 $D=0
M2083 173 94 604 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=6480 $D=0
M2084 174 94 605 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=148790 $Y=11110 $D=0
M2085 606 95 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=1850 $D=0
M2086 607 95 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=6480 $D=0
M2087 608 95 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=149170 $Y=11110 $D=0
M2088 609 603 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=1850 $D=0
M2089 610 604 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=6480 $D=0
M2090 611 605 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=149905 $Y=11110 $D=0
M2091 167 609 1023 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=1850 $D=0
M2092 173 610 1024 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=6480 $D=0
M2093 174 611 1025 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=150640 $Y=11110 $D=0
M2094 612 1023 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=1850 $D=0
M2095 613 1024 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=6480 $D=0
M2096 614 1025 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=151020 $Y=11110 $D=0
M2097 609 94 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=1850 $D=0
M2098 610 94 613 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=6480 $D=0
M2099 611 94 614 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=151465 $Y=11110 $D=0
M2100 612 606 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=1850 $D=0
M2101 613 607 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=6480 $D=0
M2102 614 608 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=152275 $Y=11110 $D=0
M2103 255 615 612 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=1850 $D=0
M2104 256 616 613 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=6480 $D=0
M2105 257 617 614 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=152795 $Y=11110 $D=0
M2106 615 96 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=1850 $D=0
M2107 616 96 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=6480 $D=0
M2108 617 96 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=153530 $Y=11110 $D=0
M2109 167 97 618 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=1850 $D=0
M2110 173 97 619 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=6480 $D=0
M2111 174 97 620 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=154190 $Y=11110 $D=0
M2112 621 98 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=1850 $D=0
M2113 622 98 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=6480 $D=0
M2114 623 98 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=154570 $Y=11110 $D=0
M2115 624 618 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=1850 $D=0
M2116 625 619 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=6480 $D=0
M2117 626 620 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=155305 $Y=11110 $D=0
M2118 167 624 1026 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=1850 $D=0
M2119 173 625 1027 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=6480 $D=0
M2120 174 626 1028 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=156040 $Y=11110 $D=0
M2121 627 1026 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=1850 $D=0
M2122 628 1027 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=6480 $D=0
M2123 629 1028 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=156420 $Y=11110 $D=0
M2124 624 97 627 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=1850 $D=0
M2125 625 97 628 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=6480 $D=0
M2126 626 97 629 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=156865 $Y=11110 $D=0
M2127 627 621 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=1850 $D=0
M2128 628 622 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=6480 $D=0
M2129 629 623 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=157675 $Y=11110 $D=0
M2130 255 630 627 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=1850 $D=0
M2131 256 631 628 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=6480 $D=0
M2132 257 632 629 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=158195 $Y=11110 $D=0
M2133 630 99 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=1850 $D=0
M2134 631 99 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=6480 $D=0
M2135 632 99 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=158930 $Y=11110 $D=0
M2136 167 100 633 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=1850 $D=0
M2137 173 100 634 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=6480 $D=0
M2138 174 100 635 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=159590 $Y=11110 $D=0
M2139 636 101 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=1850 $D=0
M2140 637 101 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=6480 $D=0
M2141 638 101 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=159970 $Y=11110 $D=0
M2142 639 633 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=1850 $D=0
M2143 640 634 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=6480 $D=0
M2144 641 635 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=160705 $Y=11110 $D=0
M2145 167 639 1029 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=1850 $D=0
M2146 173 640 1030 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=6480 $D=0
M2147 174 641 1031 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=161440 $Y=11110 $D=0
M2148 642 1029 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=1850 $D=0
M2149 643 1030 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=6480 $D=0
M2150 644 1031 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=161820 $Y=11110 $D=0
M2151 639 100 642 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=1850 $D=0
M2152 640 100 643 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=6480 $D=0
M2153 641 100 644 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=162265 $Y=11110 $D=0
M2154 642 636 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=1850 $D=0
M2155 643 637 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=6480 $D=0
M2156 644 638 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=163075 $Y=11110 $D=0
M2157 255 645 642 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=1850 $D=0
M2158 256 646 643 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=6480 $D=0
M2159 257 647 644 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=163595 $Y=11110 $D=0
M2160 645 102 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=1850 $D=0
M2161 646 102 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=6480 $D=0
M2162 647 102 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=164330 $Y=11110 $D=0
M2163 167 103 648 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=1850 $D=0
M2164 173 103 649 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=6480 $D=0
M2165 174 103 650 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=164990 $Y=11110 $D=0
M2166 651 104 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=1850 $D=0
M2167 652 104 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=6480 $D=0
M2168 653 104 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=165370 $Y=11110 $D=0
M2169 654 648 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=1850 $D=0
M2170 655 649 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=6480 $D=0
M2171 656 650 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=166105 $Y=11110 $D=0
M2172 167 654 1032 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=1850 $D=0
M2173 173 655 1033 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=6480 $D=0
M2174 174 656 1034 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=166840 $Y=11110 $D=0
M2175 657 1032 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=1850 $D=0
M2176 658 1033 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=6480 $D=0
M2177 659 1034 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=167220 $Y=11110 $D=0
M2178 654 103 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=1850 $D=0
M2179 655 103 658 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=6480 $D=0
M2180 656 103 659 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=167665 $Y=11110 $D=0
M2181 657 651 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=1850 $D=0
M2182 658 652 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=6480 $D=0
M2183 659 653 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=168475 $Y=11110 $D=0
M2184 255 660 657 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=1850 $D=0
M2185 256 661 658 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=6480 $D=0
M2186 257 662 659 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=168995 $Y=11110 $D=0
M2187 660 105 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=1850 $D=0
M2188 661 105 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=6480 $D=0
M2189 662 105 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=169730 $Y=11110 $D=0
M2190 167 106 663 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=1850 $D=0
M2191 173 106 664 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=6480 $D=0
M2192 174 106 665 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=170390 $Y=11110 $D=0
M2193 666 107 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=1850 $D=0
M2194 667 107 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=6480 $D=0
M2195 668 107 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=170770 $Y=11110 $D=0
M2196 669 663 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=1850 $D=0
M2197 670 664 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=6480 $D=0
M2198 671 665 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=171505 $Y=11110 $D=0
M2199 167 669 1035 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=1850 $D=0
M2200 173 670 1036 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=6480 $D=0
M2201 174 671 1037 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=172240 $Y=11110 $D=0
M2202 672 1035 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=1850 $D=0
M2203 673 1036 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=6480 $D=0
M2204 674 1037 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=172620 $Y=11110 $D=0
M2205 669 106 672 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=1850 $D=0
M2206 670 106 673 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=6480 $D=0
M2207 671 106 674 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=173065 $Y=11110 $D=0
M2208 672 666 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=1850 $D=0
M2209 673 667 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=6480 $D=0
M2210 674 668 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=173875 $Y=11110 $D=0
M2211 255 675 672 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=1850 $D=0
M2212 256 676 673 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=6480 $D=0
M2213 257 677 674 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=174395 $Y=11110 $D=0
M2214 675 108 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=1850 $D=0
M2215 676 108 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=6480 $D=0
M2216 677 108 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=175130 $Y=11110 $D=0
M2217 167 109 678 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=1850 $D=0
M2218 173 109 679 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=6480 $D=0
M2219 174 109 680 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=175790 $Y=11110 $D=0
M2220 681 110 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=1850 $D=0
M2221 682 110 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=6480 $D=0
M2222 683 110 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=176170 $Y=11110 $D=0
M2223 684 678 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=1850 $D=0
M2224 685 679 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=6480 $D=0
M2225 686 680 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=176905 $Y=11110 $D=0
M2226 167 684 1038 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=1850 $D=0
M2227 173 685 1039 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=6480 $D=0
M2228 174 686 1040 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=177640 $Y=11110 $D=0
M2229 687 1038 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=1850 $D=0
M2230 688 1039 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=6480 $D=0
M2231 689 1040 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=178020 $Y=11110 $D=0
M2232 684 109 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=1850 $D=0
M2233 685 109 688 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=6480 $D=0
M2234 686 109 689 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=178465 $Y=11110 $D=0
M2235 687 681 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=1850 $D=0
M2236 688 682 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=6480 $D=0
M2237 689 683 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=179275 $Y=11110 $D=0
M2238 255 690 687 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=1850 $D=0
M2239 256 691 688 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=6480 $D=0
M2240 257 692 689 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=179795 $Y=11110 $D=0
M2241 690 113 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=1850 $D=0
M2242 691 113 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=6480 $D=0
M2243 692 113 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=180530 $Y=11110 $D=0
M2244 167 114 693 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=1850 $D=0
M2245 173 114 694 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=6480 $D=0
M2246 174 114 695 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=181190 $Y=11110 $D=0
M2247 696 115 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=1850 $D=0
M2248 697 115 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=6480 $D=0
M2249 698 115 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=181570 $Y=11110 $D=0
M2250 699 693 234 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=1850 $D=0
M2251 700 694 235 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=6480 $D=0
M2252 701 695 236 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=182305 $Y=11110 $D=0
M2253 167 699 1041 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=1850 $D=0
M2254 173 700 1042 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=6480 $D=0
M2255 174 701 1043 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=183040 $Y=11110 $D=0
M2256 702 1041 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=1850 $D=0
M2257 703 1042 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=6480 $D=0
M2258 704 1043 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=183420 $Y=11110 $D=0
M2259 699 114 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=1850 $D=0
M2260 700 114 703 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=6480 $D=0
M2261 701 114 704 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=183865 $Y=11110 $D=0
M2262 702 696 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=1850 $D=0
M2263 703 697 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=6480 $D=0
M2264 704 698 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=184675 $Y=11110 $D=0
M2265 255 705 702 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=1850 $D=0
M2266 256 706 703 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=6480 $D=0
M2267 257 707 704 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=185195 $Y=11110 $D=0
M2268 705 118 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=1850 $D=0
M2269 706 118 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=6480 $D=0
M2270 707 118 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=185930 $Y=11110 $D=0
M2271 167 119 708 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=1850 $D=0
M2272 173 119 709 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=6480 $D=0
M2273 174 119 710 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=186590 $Y=11110 $D=0
M2274 711 120 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=1850 $D=0
M2275 712 120 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=6480 $D=0
M2276 713 120 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=186970 $Y=11110 $D=0
M2277 7 711 249 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=1850 $D=0
M2278 8 712 250 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=6480 $D=0
M2279 9 713 251 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=187705 $Y=11110 $D=0
M2280 255 708 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=1850 $D=0
M2281 256 709 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=6480 $D=0
M2282 257 710 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=188225 $Y=11110 $D=0
M2283 167 717 714 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=1850 $D=0
M2284 173 718 715 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=6480 $D=0
M2285 174 719 716 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=188960 $Y=11110 $D=0
M2286 717 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=1850 $D=0
M2287 718 121 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=6480 $D=0
M2288 719 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=189340 $Y=11110 $D=0
M2289 1044 249 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=1850 $D=0
M2290 1045 250 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=6480 $D=0
M2291 1046 251 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=190000 $Y=11110 $D=0
M2292 720 717 1044 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=1850 $D=0
M2293 721 718 1045 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=6480 $D=0
M2294 722 719 1046 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=190445 $Y=11110 $D=0
M2295 167 720 122 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=1850 $D=0
M2296 173 721 723 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=6480 $D=0
M2297 174 722 724 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=191180 $Y=11110 $D=0
M2298 1047 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=1850 $D=0
M2299 1048 723 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=6480 $D=0
M2300 1049 724 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=191560 $Y=11110 $D=0
M2301 720 714 1047 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=1850 $D=0
M2302 721 715 1048 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=6480 $D=0
M2303 722 716 1049 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=192280 $Y=11110 $D=0
M2304 167 728 725 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=1850 $D=0
M2305 173 729 726 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=6480 $D=0
M2306 174 730 727 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=192955 $Y=11110 $D=0
M2307 728 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=1850 $D=0
M2308 729 121 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=6480 $D=0
M2309 730 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=193335 $Y=11110 $D=0
M2310 1050 255 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=1850 $D=0
M2311 1051 256 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=6480 $D=0
M2312 1052 257 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=193995 $Y=11110 $D=0
M2313 731 728 1050 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=1850 $D=0
M2314 732 729 1051 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=6480 $D=0
M2315 733 730 1052 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=194440 $Y=11110 $D=0
M2316 167 731 123 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=1850 $D=0
M2317 173 732 124 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=6480 $D=0
M2318 174 733 125 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=195175 $Y=11110 $D=0
M2319 1053 123 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=1850 $D=0
M2320 1054 124 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=6480 $D=0
M2321 1055 125 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=195555 $Y=11110 $D=0
M2322 731 725 1053 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=1850 $D=0
M2323 732 726 1054 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=6480 $D=0
M2324 733 727 1055 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=196275 $Y=11110 $D=0
M2325 734 126 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=1850 $D=0
M2326 735 126 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=6480 $D=0
M2327 736 126 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=196950 $Y=11110 $D=0
M2328 737 126 122 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=1850 $D=0
M2329 738 126 723 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=6480 $D=0
M2330 739 126 724 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=197685 $Y=11110 $D=0
M2331 127 734 737 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=1850 $D=0
M2332 128 735 738 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=6480 $D=0
M2333 129 736 739 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=198205 $Y=11110 $D=0
M2334 740 130 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=1850 $D=0
M2335 741 130 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=6480 $D=0
M2336 742 130 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=198945 $Y=11110 $D=0
M2337 743 130 123 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=1850 $D=0
M2338 744 130 124 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=6480 $D=0
M2339 745 130 125 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=199680 $Y=11110 $D=0
M2340 1056 740 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=1850 $D=0
M2341 1057 741 744 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=6480 $D=0
M2342 1058 742 745 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.78e-14 PD=7.05e-07 PS=7.8e-07 $X=200200 $Y=11110 $D=0
M2343 167 123 1056 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=1850 $D=0
M2344 173 124 1057 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=6480 $D=0
M2345 174 125 1058 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=3.105e-14 PD=5.6e-07 PS=7.05e-07 $X=200645 $Y=11110 $D=0
M2346 746 131 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=1850 $D=0
M2347 747 131 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=6480 $D=0
M2348 748 131 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=201305 $Y=11110 $D=0
M2349 749 131 743 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=1850 $D=0
M2350 750 131 744 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=6480 $D=0
M2351 751 131 745 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=202040 $Y=11110 $D=0
M2352 14 746 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=1850 $D=0
M2353 15 747 750 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=6480 $D=0
M2354 16 748 751 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=202560 $Y=11110 $D=0
M2355 755 752 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=1850 $D=0
M2356 756 753 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=6480 $D=0
M2357 757 754 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=203300 $Y=11110 $D=0
M2358 167 761 758 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=1850 $D=0
M2359 173 762 759 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=6480 $D=0
M2360 174 763 760 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=203960 $Y=11110 $D=0
M2361 764 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=1850 $D=0
M2362 765 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=6480 $D=0
M2363 766 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=204340 $Y=11110 $D=0
M2364 761 737 752 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=1850 $D=0
M2365 762 738 753 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=6480 $D=0
M2366 763 739 754 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=205075 $Y=11110 $D=0
M2367 755 764 761 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=1850 $D=0
M2368 756 765 762 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=6480 $D=0
M2369 757 766 763 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=205595 $Y=11110 $D=0
M2370 767 758 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=1850 $D=0
M2371 768 759 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=6480 $D=0
M2372 769 760 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=206330 $Y=11110 $D=0
M2373 770 758 749 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=1850 $D=0
M2374 771 759 750 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=6480 $D=0
M2375 772 760 751 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=207065 $Y=11110 $D=0
M2376 737 767 770 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=1850 $D=0
M2377 738 768 771 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=6480 $D=0
M2378 739 769 772 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=207585 $Y=11110 $D=0
M2379 773 770 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=1850 $D=0
M2380 774 771 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=6480 $D=0
M2381 775 772 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208320 $Y=11110 $D=0
M2382 776 758 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=1850 $D=0
M2383 777 759 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=6480 $D=0
M2384 778 760 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=208980 $Y=11110 $D=0
M2385 779 758 773 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=1850 $D=0
M2386 780 759 774 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=6480 $D=0
M2387 781 760 775 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=209715 $Y=11110 $D=0
M2388 749 776 779 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=1850 $D=0
M2389 750 777 780 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=6480 $D=0
M2390 751 778 781 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=210235 $Y=11110 $D=0
M2391 1074 737 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=1490 $D=0
M2392 1075 738 173 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=6120 $D=0
M2393 1076 739 174 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=210970 $Y=10750 $D=0
M2394 782 749 1074 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=1490 $D=0
M2395 783 750 1075 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=6120 $D=0
M2396 784 751 1076 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=211350 $Y=10750 $D=0
M2397 785 779 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=1850 $D=0
M2398 786 780 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=6480 $D=0
M2399 787 781 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=212010 $Y=11110 $D=0
M2400 788 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=1850 $D=0
M2401 789 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=6480 $D=0
M2402 790 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=212670 $Y=11110 $D=0
M2403 167 749 788 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=1850 $D=0
M2404 173 750 789 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=6480 $D=0
M2405 174 751 790 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=213050 $Y=11110 $D=0
M2406 791 737 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=1850 $D=0
M2407 792 738 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=6480 $D=0
M2408 793 739 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=213710 $Y=11110 $D=0
M2409 167 749 791 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=1850 $D=0
M2410 173 750 792 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=6480 $D=0
M2411 174 751 793 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=214090 $Y=11110 $D=0
M2412 1077 737 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=1670 $D=0
M2413 1078 738 173 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=6300 $D=0
M2414 1079 739 174 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=214750 $Y=10930 $D=0
M2415 797 749 1077 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=1670 $D=0
M2416 798 750 1078 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=6300 $D=0
M2417 799 751 1079 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=215130 $Y=10930 $D=0
M2418 167 791 797 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=1850 $D=0
M2419 173 792 798 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=6480 $D=0
M2420 174 793 799 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.845e-14 AS=3.735e-14 PD=5.65e-07 PS=8.55e-07 $X=215545 $Y=11110 $D=0
M2421 800 135 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=1850 $D=0
M2422 801 135 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=6480 $D=0
M2423 802 135 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=216210 $Y=11110 $D=0
M2424 803 135 782 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=1850 $D=0
M2425 804 135 783 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=6480 $D=0
M2426 805 135 784 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=216945 $Y=11110 $D=0
M2427 788 800 803 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=1850 $D=0
M2428 789 801 804 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=6480 $D=0
M2429 790 802 805 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=217465 $Y=11110 $D=0
M2430 806 135 785 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=1850 $D=0
M2431 807 135 786 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=6480 $D=0
M2432 808 135 787 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=218275 $Y=11110 $D=0
M2433 797 800 806 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=1850 $D=0
M2434 798 801 807 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=6480 $D=0
M2435 799 802 808 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=218795 $Y=11110 $D=0
M2436 809 136 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=1850 $D=0
M2437 810 136 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=6480 $D=0
M2438 811 136 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=219530 $Y=11110 $D=0
M2439 812 136 806 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=1850 $D=0
M2440 813 136 807 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=6480 $D=0
M2441 814 136 808 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=220265 $Y=11110 $D=0
M2442 803 809 812 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=1850 $D=0
M2443 804 810 813 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=6480 $D=0
M2444 805 811 814 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=220785 $Y=11110 $D=0
M2445 17 812 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=1850 $D=0
M2446 18 813 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=6480 $D=0
M2447 19 814 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=221520 $Y=11110 $D=0
M2448 815 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=1850 $D=0
M2449 816 137 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=6480 $D=0
M2450 817 137 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=222180 $Y=11110 $D=0
M2451 818 137 138 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=1850 $D=0
M2452 819 137 139 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=6480 $D=0
M2453 820 137 140 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=222915 $Y=11110 $D=0
M2454 141 815 818 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=1850 $D=0
M2455 142 816 819 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=6480 $D=0
M2456 138 817 820 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=223435 $Y=11110 $D=0
M2457 821 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=1850 $D=0
M2458 822 137 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=6480 $D=0
M2459 823 137 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=224170 $Y=11110 $D=0
M2460 824 137 143 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=1850 $D=0
M2461 825 137 144 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=6480 $D=0
M2462 826 137 145 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=224905 $Y=11110 $D=0
M2463 141 821 824 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=1850 $D=0
M2464 141 822 825 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=6480 $D=0
M2465 146 823 826 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=225425 $Y=11110 $D=0
M2466 827 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=1850 $D=0
M2467 828 137 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=6480 $D=0
M2468 829 137 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=226160 $Y=11110 $D=0
M2469 830 137 134 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=1850 $D=0
M2470 831 137 133 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=6480 $D=0
M2471 832 137 132 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=226895 $Y=11110 $D=0
M2472 141 827 830 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=1850 $D=0
M2473 141 828 831 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=6480 $D=0
M2474 141 829 832 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=227415 $Y=11110 $D=0
M2475 833 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=1850 $D=0
M2476 834 137 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=6480 $D=0
M2477 835 137 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=228150 $Y=11110 $D=0
M2478 836 137 147 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=1850 $D=0
M2479 837 137 148 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=6480 $D=0
M2480 838 137 149 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=228885 $Y=11110 $D=0
M2481 141 833 836 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=1850 $D=0
M2482 141 834 837 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=6480 $D=0
M2483 141 835 838 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=229405 $Y=11110 $D=0
M2484 839 137 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=1850 $D=0
M2485 840 137 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=6480 $D=0
M2486 841 137 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=230140 $Y=11110 $D=0
M2487 842 137 150 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=1850 $D=0
M2488 843 137 151 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=6480 $D=0
M2489 844 137 152 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=230875 $Y=11110 $D=0
M2490 141 839 842 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=1850 $D=0
M2491 141 840 843 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=6480 $D=0
M2492 141 841 844 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=231395 $Y=11110 $D=0
M2493 167 737 1059 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=1850 $D=0
M2494 173 738 1060 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=6480 $D=0
M2495 174 739 1061 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=232130 $Y=11110 $D=0
M2496 142 1059 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=1850 $D=0
M2497 138 1060 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=6480 $D=0
M2498 139 1061 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=232510 $Y=11110 $D=0
M2499 845 153 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=1850 $D=0
M2500 846 153 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=6480 $D=0
M2501 847 153 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=233170 $Y=11110 $D=0
M2502 146 153 142 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=1850 $D=0
M2503 154 153 138 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=6480 $D=0
M2504 143 153 139 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=233905 $Y=11110 $D=0
M2505 818 845 146 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=1850 $D=0
M2506 819 846 154 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=6480 $D=0
M2507 820 847 143 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=234425 $Y=11110 $D=0
M2508 848 155 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=1850 $D=0
M2509 849 155 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=6480 $D=0
M2510 850 155 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=235160 $Y=11110 $D=0
M2511 156 155 146 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=1850 $D=0
M2512 157 155 154 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=6480 $D=0
M2513 158 155 143 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=235895 $Y=11110 $D=0
M2514 824 848 156 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=1850 $D=0
M2515 825 849 157 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=6480 $D=0
M2516 826 850 158 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=236415 $Y=11110 $D=0
M2517 851 159 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=1850 $D=0
M2518 852 159 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=6480 $D=0
M2519 853 159 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=237150 $Y=11110 $D=0
M2520 112 159 156 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=1850 $D=0
M2521 116 159 157 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=6480 $D=0
M2522 111 159 158 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=237885 $Y=11110 $D=0
M2523 830 851 112 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=1850 $D=0
M2524 831 852 116 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=6480 $D=0
M2525 832 853 111 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=238405 $Y=11110 $D=0
M2526 854 160 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=1850 $D=0
M2527 855 160 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=6480 $D=0
M2528 856 160 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=239140 $Y=11110 $D=0
M2529 161 160 112 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=1850 $D=0
M2530 162 160 116 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=6480 $D=0
M2531 163 160 111 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=239875 $Y=11110 $D=0
M2532 836 854 161 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=1850 $D=0
M2533 837 855 162 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=6480 $D=0
M2534 838 856 163 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=240395 $Y=11110 $D=0
M2535 857 164 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=1850 $D=0
M2536 858 164 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=6480 $D=0
M2537 859 164 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=241130 $Y=11110 $D=0
M2538 213 164 161 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=1850 $D=0
M2539 214 164 162 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=6480 $D=0
M2540 215 164 163 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=241865 $Y=11110 $D=0
M2541 842 857 213 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=1850 $D=0
M2542 843 858 214 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=6480 $D=0
M2543 844 859 215 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=242385 $Y=11110 $D=0
M2544 860 165 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=1850 $D=0
M2545 861 165 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=6480 $D=0
M2546 862 165 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=243120 $Y=11110 $D=0
M2547 166 165 123 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=1850 $D=0
M2548 863 165 124 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=6480 $D=0
M2549 864 165 125 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=243855 $Y=11110 $D=0
M2550 14 860 166 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=1850 $D=0
M2551 15 861 863 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=6480 $D=0
M2552 16 862 864 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=244375 $Y=11110 $D=0
M2553 865 122 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=1850 $D=0
M2554 866 723 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=6480 $D=0
M2555 867 724 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=245110 $Y=11110 $D=0
M2556 167 166 865 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=1850 $D=0
M2557 173 863 866 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=6480 $D=0
M2558 174 864 867 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=245490 $Y=11110 $D=0
M2559 1080 122 167 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=1670 $D=0
M2560 1081 723 173 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=6300 $D=0
M2561 1082 724 174 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.7e-14 PD=8.2e-07 PS=7.4e-07 $X=246150 $Y=10930 $D=0
M2562 871 166 1080 167 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=1670 $D=0
M2563 872 863 1081 173 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=6300 $D=0
M2564 873 864 1082 174 PMOS_VTL L=5e-08 W=2.7e-07 AD=3.735e-14 AS=3.78e-14 PD=8.55e-07 PS=8.2e-07 $X=246530 $Y=10930 $D=0
M2565 167 865 871 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=1850 $D=0
M2566 173 866 872 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=6480 $D=0
M2567 174 867 873 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.835e-14 AS=3.735e-14 PD=6.75e-07 PS=8.55e-07 $X=246945 $Y=11110 $D=0
M2568 1062 167 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=1850 $D=0
M2569 1063 874 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=6480 $D=0
M2570 1064 875 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.835e-14 PD=6.4e-07 PS=6.75e-07 $X=247360 $Y=11110 $D=0
M2571 167 871 1062 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=1850 $D=0
M2572 173 872 1063 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=6480 $D=0
M2573 174 873 1064 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=247740 $Y=11110 $D=0
M2574 874 1062 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=1850 $D=0
M2575 875 1063 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=6480 $D=0
M2576 168 1064 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=248400 $Y=11110 $D=0
M2577 1083 122 167 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=1490 $D=0
M2578 1084 723 173 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=6120 $D=0
M2579 1085 724 174 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.6e-14 PD=1e-06 PS=9.2e-07 $X=249060 $Y=10750 $D=0
M2580 876 879 1083 167 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=1490 $D=0
M2581 877 880 1084 173 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=6120 $D=0
M2582 878 881 1085 174 PMOS_VTL L=5e-08 W=3.6e-07 AD=3.6e-14 AS=5.04e-14 PD=9.2e-07 PS=1e-06 $X=249440 $Y=10750 $D=0
M2583 879 166 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=1850 $D=0
M2584 880 863 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=6480 $D=0
M2585 881 864 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=250100 $Y=11110 $D=0
M2586 882 876 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=1850 $D=0
M2587 883 877 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=6480 $D=0
M2588 884 878 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=250760 $Y=11110 $D=0
M2589 167 167 882 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=1850 $D=0
M2590 173 874 883 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=6480 $D=0
M2591 174 875 884 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=251140 $Y=11110 $D=0
M2592 887 7 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=1850 $D=0
M2593 888 885 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=6480 $D=0
M2594 889 886 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=251800 $Y=11110 $D=0
M2595 885 882 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=1850 $D=0
M2596 886 883 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=6480 $D=0
M2597 169 884 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=252460 $Y=11110 $D=0
M2598 167 887 885 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=1850 $D=0
M2599 173 888 886 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=6480 $D=0
M2600 174 889 169 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=252840 $Y=11110 $D=0
M2601 892 890 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=1850 $D=0
M2602 893 891 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=6480 $D=0
M2603 894 170 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=253500 $Y=11110 $D=0
M2604 167 898 895 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=1850 $D=0
M2605 173 899 896 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=6480 $D=0
M2606 174 900 897 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=254160 $Y=11110 $D=0
M2607 901 127 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=1850 $D=0
M2608 902 128 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=6480 $D=0
M2609 903 129 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=254540 $Y=11110 $D=0
M2610 898 127 890 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=1850 $D=0
M2611 899 128 891 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=6480 $D=0
M2612 900 129 170 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=255275 $Y=11110 $D=0
M2613 892 901 898 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=1850 $D=0
M2614 893 902 899 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=6480 $D=0
M2615 894 903 900 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=255795 $Y=11110 $D=0
M2616 904 895 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=1850 $D=0
M2617 905 896 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=6480 $D=0
M2618 906 897 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=256530 $Y=11110 $D=0
M2619 907 895 7 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=1850 $D=0
M2620 890 896 8 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=6480 $D=0
M2621 891 897 9 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=257265 $Y=11110 $D=0
M2622 127 904 907 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=1850 $D=0
M2623 128 905 890 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=6480 $D=0
M2624 129 906 891 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=257785 $Y=11110 $D=0
M2625 908 907 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=1850 $D=0
M2626 909 890 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=6480 $D=0
M2627 910 891 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=258520 $Y=11110 $D=0
M2628 911 895 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=1850 $D=0
M2629 912 896 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=6480 $D=0
M2630 913 897 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=259180 $Y=11110 $D=0
M2631 216 895 908 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=1850 $D=0
M2632 217 896 909 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=6480 $D=0
M2633 218 897 910 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=259915 $Y=11110 $D=0
M2634 7 911 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=1850 $D=0
M2635 8 912 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=6480 $D=0
M2636 9 913 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=260435 $Y=11110 $D=0
M2637 914 171 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=1850 $D=0
M2638 915 171 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=6480 $D=0
M2639 916 171 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=261170 $Y=11110 $D=0
M2640 917 171 216 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=1850 $D=0
M2641 918 171 217 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=6480 $D=0
M2642 919 171 218 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=261905 $Y=11110 $D=0
M2643 17 914 917 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=1850 $D=0
M2644 18 915 918 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=6480 $D=0
M2645 19 916 919 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=262425 $Y=11110 $D=0
M2646 920 172 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=1850 $D=0
M2647 921 172 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=6480 $D=0
M2648 922 172 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=263160 $Y=11110 $D=0
M2649 923 172 917 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=1850 $D=0
M2650 172 172 918 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=6480 $D=0
M2651 172 172 919 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=263895 $Y=11110 $D=0
M2652 7 920 923 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=1850 $D=0
M2653 173 921 172 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=6480 $D=0
M2654 174 922 172 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=264415 $Y=11110 $D=0
M2655 924 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=1850 $D=0
M2656 925 121 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=6480 $D=0
M2657 926 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=265150 $Y=11110 $D=0
M2658 167 924 927 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=1850 $D=0
M2659 173 925 928 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=6480 $D=0
M2660 174 926 929 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=265810 $Y=11110 $D=0
M2661 930 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=1850 $D=0
M2662 931 121 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=6480 $D=0
M2663 932 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=266190 $Y=11110 $D=0
M2664 933 927 923 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=1850 $D=0
M2665 934 928 172 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=6480 $D=0
M2666 935 929 172 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=266925 $Y=11110 $D=0
M2667 167 933 1065 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=1850 $D=0
M2668 173 934 1066 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=6480 $D=0
M2669 174 935 1067 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=267660 $Y=11110 $D=0
M2670 936 1065 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=1850 $D=0
M2671 937 1066 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=6480 $D=0
M2672 938 1067 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=268040 $Y=11110 $D=0
M2673 933 924 936 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=1850 $D=0
M2674 934 925 937 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=6480 $D=0
M2675 935 926 938 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=268485 $Y=11110 $D=0
M2676 939 930 936 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=1850 $D=0
M2677 940 931 937 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=6480 $D=0
M2678 941 932 938 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=269295 $Y=11110 $D=0
M2679 167 945 942 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=1850 $D=0
M2680 173 946 943 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=6480 $D=0
M2681 174 947 944 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=270030 $Y=11110 $D=0
M2682 945 121 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=1850 $D=0
M2683 946 121 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=6480 $D=0
M2684 947 121 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=270410 $Y=11110 $D=0
M2685 1068 939 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=1850 $D=0
M2686 1069 940 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=6480 $D=0
M2687 1070 941 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=271070 $Y=11110 $D=0
M2688 948 945 1068 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=1850 $D=0
M2689 949 946 1069 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=6480 $D=0
M2690 950 947 1070 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=271515 $Y=11110 $D=0
M2691 167 948 127 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=1850 $D=0
M2692 173 949 128 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=6480 $D=0
M2693 174 950 129 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=272250 $Y=11110 $D=0
M2694 1071 127 167 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=1850 $D=0
M2695 1072 128 173 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=6480 $D=0
M2696 1073 129 174 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=272630 $Y=11110 $D=0
M2697 948 942 1071 167 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=1850 $D=0
M2698 949 943 1072 173 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=6480 $D=0
M2699 950 944 1073 174 PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=273350 $Y=11110 $D=0
.ENDS
***************************************
.SUBCKT datapath 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 vdd! 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 vss! 60
+ 61 62 63 64 shift_out<8> shift_out<18> shift_out<28> shift_out<38> shift_out<48> shift_out<9> shift_out<114> mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> cmp_out imm<2>
+ imm<1> imm<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26>
+ rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20>
+ rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13>
+ rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6>
+ rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk
+ dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel alu_inv_rs2 alu_mux_2_sel alu_cin shift_out<13> shift_out<3> shift_out<2> shift_out<7> shift_out<12> alu_op<0> alu_op<1> shift_out<16> dmem_addr<2> dmem_addr<1> dmem_addr<0> shift_dir shift_out<10>
+ shift_out<5> shift_out<0> shift_out<15> shift_out<6> shift_out<1> shift_out<21> shift_out<11> 213 shift_out<27> shift_out<22> shift_out<53> shift_out<43> shift_out<94> shift_out<89> shift_out<84> shift_amount<0> shift_amount<1> shift_amount<2> shift_amount<3> shift_amount<4>
+ shift_out<14> shift_out<4> cmp_mux_sel cmp_eq cmp_lt pc_mux_sel rst imem_addr<2> imem_addr<1> imem_addr<0> dmem_rdata<4> dmem_rdata<3> imm<4> imm<3> dmem_wdata<4> dmem_wdata<3> shift_out<23> shift_out<17> 248 shift_out<26>
+ dmem_addr<3> dmem_addr<4> shift_out<20> shift_out<25> shift_out<31> 255 shift_out<63> shift_out<58> shift_out<104> shift_out<99> shift_out<24> shift_out<19> imem_addr<4> imem_addr<3> dmem_rdata<6> dmem_rdata<5> imm<6> imm<5> dmem_wdata<6> dmem_wdata<5>
+ shift_out<33> shift_out<32> shift_out<36> dmem_addr<6> dmem_addr<5> shift_out<30> shift_out<35> shift_out<41> shift_out<52> shift_out<47> shift_out<73> shift_out<68> shift_out<109> imem_addr<10> shift_out<29> imem_addr<6> imem_addr<5> dmem_rdata<8> dmem_rdata<7> imm<8>
+ imm<7> dmem_wdata<8> dmem_wdata<7> shift_out<62> shift_out<83> shift_out<57> shift_out<42> shift_out<37> shift_out<46> dmem_addr<8> dmem_addr<7> shift_out<40> shift_out<45> shift_out<51> shift_out<78> shift_out<124> shift_out<119> shift_out<44> shift_out<39> dmem_rdata<10>
+ dmem_rdata<9> imm<10> imm<9> dmem_wdata<10> dmem_wdata<9> shift_out<92> shift_out<72> shift_out<87> shift_out<67> dmem_addr<9> dmem_addr<10> shift_out<50> shift_out<55> shift_out<61> shift_out<134> shift_out<129> shift_out<54> shift_out<49> dmem_rdata<12> dmem_rdata<11>
+ imm<12> imm<11> dmem_wdata<12> dmem_wdata<11> shift_out<82> shift_out<102> shift_out<77> shift_out98> dmem_addr<11> dmem_addr<12> shift_out<60> shift_out<65> shift_out<71> shift_out<144> shift_out<139> shift_out<64> shift_out<59> dmem_rdata<14> dmem_rdata<13> imm<14>
+ imm<13> shift_out<112> shift_out<107> dmem_wdata<14> dmem_wdata<13> dmem_addr<14> dmem_addr<13> shift_out<70> shift_out<75> shift_out<81> shift_out<154> shift_out<149> shift_out<74> shift_out<69> dmem_rdata<16> dmem_rdata<15> imm<16> imm<15> shift_out<123> shift_out<117>
+ dmem_wdata<16> dmem_wdata<15> shift_out<86> dmem_addr<16> dmem_addr<15> shift_out<80> shift_out<91> shift_msb shift_out<159> shift_out<85> shift_out<79> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> imm<20> imm<19> imm<18> imm<17> shift_out<138>
+ shift_out<133> shift_out<128> dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> shift_out<96> shift_out<106> dmem_addr<17> dmem_addr<20> dmem_addr<19> dmem_addr<18> shift_out<95> shift_out<90> shift_out<105> shift_out<100> shift_out<111> shift_out<101> shift_out<122> shift_out<143>
+ dmem_rdata<22> dmem_rdata<21> imm<22> imm<21> shift_out<127> shift_out<148> dmem_wdata<22> dmem_wdata<21> 450 shift_out<116> dmem_addr<22> dmem_addr<21> shift_out<115> shift_out<110> shift_out<121> shift_out<132> shift_out<153> imem_addr<22> dmem_rdata<24> dmem_rdata<23>
+ imm<24> imm<23> shift_out<137> shift_out<158> dmem_wdata<24> dmem_wdata<23> shift_out<126> dmem_addr<24> dmem_addr<23> shift_out<125> shift_out<120> shift_out<131> shift_out<142> imem_addr<24> imem_addr<23> dmem_rdata<26> dmem_rdata<25> imm<26> imm<25> dmem_wdata<26>
+ dmem_wdata<25> shift_out<136> dmem_addr<26> dmem_addr<25> shift_out<135> shift_out<130> shift_out<141> shift_out<152> shift_out<147> imem_addr<26> imem_addr<25> dmem_rdata<28> dmem_rdata<27> imm<28> imm<27> dmem_wdata<28> dmem_wdata<27> shift_out<146> dmem_addr<28> dmem_addr<27>
+ shift_out<145> shift_out<140> shift_out<151> shift_out<157> imem_addr<28> imem_addr<27> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> imm<31> imm<30> imm<29> dmem_wdata<31> dmem_wdata<30> dmem_wdata<29> dmem_addr<31> dmem_addr<30> dmem_addr<29> shift_out<150> shift_out<155>
+ shift_out<156> cmp_a_31 cmp_b_31 imem_addr<31> imem_addr<30> imem_addr<29>
** N=538 EP=486 IP=2688 FDC=28800
X0 mem_mux_sel<0> dmem_rdata<2> dmem_rdata<1> dmem_rdata<0> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 1 3 cmp_out imm<2> imm<1> imm<0> dmem_addr<2> dmem_addr<1> dmem_addr<0> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31>
+ rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24>
+ rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18>
+ rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11>
+ rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4>
+ rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<2> dmem_wdata<1> dmem_wdata<0> alu_mux_1_sel imem_addr<2> imem_addr<1>
+ imem_addr<0> alu_inv_rs2 alu_mux_2_sel shift_amount<2> shift_amount<1> shift_amount<0> alu_cin 191 shift_out<13> shift_out<8> shift_out<3> shift_out<2> shift_out<7> shift_out<12> alu_op<0> alu_op<1> shift_dir shift_out<5> shift_out<0> 5
+ shift_out<15> shift_out<10> shift_out<1> shift_out<21> shift_out<16> shift_out<11> 213 shift_out<27> shift_out<22> shift_out<53> shift_out<48> shift_out<43> shift_out<94> shift_out<89> shift_out<84> shift_out<6> shift_amount<3> shift_out<14> shift_out<9> shift_out<4>
+ shift_amount<4> cmp_mux_sel 229 cmp_eq 231 cmp_lt 2 233 pc_mux_sel rst 4 6
+ ICV_24 $T=0 0 0 0 $X=0 $Y=132400
X1 mem_mux_sel<0> dmem_rdata<4> dmem_rdata<3> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 7 9 imm<4> imm<3> dmem_addr<4> dmem_addr<3> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<4> dmem_wdata<3> alu_mux_1_sel imem_addr<4> imem_addr<3> alu_inv_rs2 alu_mux_2_sel shift_amount<4> shift_amount<3> 191
+ shift_out<23> shift_out<18> shift_out<2> shift_out<17> alu_op<0> alu_op<1> 248 shift_dir shift_out<15> shift_out<10> shift_out<25> shift_out<20> shift_out<11> shift_out<6> shift_out<31> shift_out<26> shift_out<53> 255 shift_out<63> shift_out<58>
+ shift_out<104> shift_out<99> shift_amount<0> shift_out<21> shift_out<16> shift_amount<1> shift_out<22> shift_amount<2> shift_out<24> shift_out<19> cmp_mux_sel 262 229 263 231 233 264 pc_mux_sel rst 8
+ 10
+ ICV_25 $T=0 0 0 0 $X=0 $Y=123200
X2 mem_mux_sel<0> dmem_rdata<6> dmem_rdata<5> mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 11 13 imm<6> imm<5> dmem_addr<6> dmem_addr<5> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<6> dmem_wdata<5> alu_mux_1_sel imem_addr<6> imem_addr<5> alu_inv_rs2 alu_mux_2_sel 245 shift_out<33> shift_out<28>
+ 273 shift_out<12> alu_op<0> alu_op<1> shift_dir shift_out<25> shift_out<20> shift_out<35> shift_out<30> shift_out<21> shift_out<16> shift_out<41> shift_out<36> shift_out<7> shift_out<53> shift_out<52> shift_out<47> shift_out<73> shift_out<68> shift_out<114>
+ shift_out<109> shift_amount<0> shift_out<31> shift_out<26> shift_amount<1> shift_out<32> shift_out<27> shift_amount<2> shift_amount<3> imem_addr<10> shift_out<29> shift_amount<4> cmp_mux_sel 289 262 290 263 264 291 pc_mux_sel
+ rst 12 14
+ ICV_26 $T=0 0 0 0 $X=0 $Y=114000
X3 mem_mux_sel<0> dmem_rdata<8> dmem_rdata<7> 15 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> 17 imm<8> imm<7> dmem_addr<8> dmem_addr<7> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30>
+ rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23>
+ rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16>
+ rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10>
+ rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3>
+ rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<8> dmem_wdata<7> alu_mux_1_sel imem_addr<10> alu_inv_rs2 shift_out<62> alu_mux_2_sel shift_out<83> 273 shift_out<43>
+ shift_out<38> shift_out<57> shift_out<42> alu_op<0> alu_op<1> shift_dir shift_out<35> shift_out<30> shift_out<45> shift_out<40> shift_out<31> shift_out<26> shift_out<51> shift_out<46> shift_out<22> shift_out<17> shift_out<53> shift_out<3> shift_out<78> shift_out<124>
+ shift_out<119> shift_amount<0> shift_out<41> shift_out<36> shift_amount<1> shift_out<37> shift_amount<2> shift_amount<3> shift_out<44> shift_out<39> shift_amount<4> cmp_mux_sel 317 289 318 290 291 319 pc_mux_sel rst
+ 16 18
+ ICV_27 $T=0 0 0 0 $X=0 $Y=104600
X4 mem_mux_sel<0> dmem_rdata<10> dmem_rdata<9> dmem_rdata<7> 19 21 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<10> imm<9> dmem_addr<10> dmem_addr<9> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<10> dmem_wdata<9> shift_out<92> alu_mux_1_sel shift_out<72> imem_addr<10> alu_inv_rs2 shift_out<87> shift_out<67>
+ alu_mux_2_sel 302 shift_out<53> shift_out<48> 330 shift_out<47> alu_op<0> alu_op<1> shift_dir shift_out<45> shift_out<40> shift_out<55> shift_out<50> shift_out<41> shift_out<36> shift_out<61> shift_out<32> shift_out<27> shift_out<13> shift_out<8>
+ shift_out<134> shift_out<129> shift_amount<0> shift_out<51> shift_out<46> shift_amount<1> shift_out<52> shift_amount<2> shift_amount<3> shift_out<54> shift_out<49> shift_amount<4> cmp_mux_sel 340 317 341 318 319 342 pc_mux_sel
+ rst 20 22
+ ICV_28 $T=0 0 0 0 $X=0 $Y=95400
X5 mem_mux_sel<0> dmem_rdata<12> dmem_rdata<11> dmem_rdata<7> 23 25 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<12> imm<11> dmem_addr<12> dmem_addr<11> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<12> dmem_wdata<11> shift_out<82> shift_out<102> shift_out<77> shift_out98> alu_mux_1_sel imem_addr<10> alu_inv_rs2
+ shift_out<62> alu_mux_2_sel 330 shift_out<63> shift_out<58> alu_op<0> alu_op<1> shift_dir shift_out<55> shift_out<50> shift_out<65> shift_out<60> shift_out<51> shift_out<46> shift_out<71> shift_out<42> shift_out<37> shift_out<23> shift_out<18> shift_out<144>
+ shift_out<139> shift_amount<0> shift_out<61> shift_out<32> shift_amount<1> shift_out<57> shift_amount<2> shift_amount<3> shift_out<64> shift_out<59> shift_amount<4> cmp_mux_sel 363 340 364 341 342 365 pc_mux_sel rst
+ vdd! 26
+ ICV_29 $T=0 0 0 0 $X=0 $Y=86200
X6 mem_mux_sel<0> dmem_rdata<14> dmem_rdata<13> dmem_rdata<7> 27 29 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<14> imm<13> dmem_addr<14> dmem_addr<13> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk shift_out<73> shift_out<92> shift_out<112> shift_out<87> shift_out<107> dmem_wdata<14> dmem_wdata<13> alu_mux_1_sel shift_out<72>
+ imem_addr<10> alu_inv_rs2 shift_out<67> alu_mux_2_sel 353 shift_out<68> 374 alu_op<0> alu_op<1> shift_dir shift_out<65> shift_out<60> shift_out<75> shift_out<70> shift_out<61> shift_out<32> shift_out<81> shift_out<52> shift_out<47> shift_out<33>
+ shift_out<28> shift_out<154> shift_out<149> shift_amount<0> shift_out<71> shift_out<42> shift_amount<1> shift_amount<2> shift_amount<3> shift_out<74> shift_out<69> shift_amount<4> cmp_mux_sel 384 363 385 364 365 386 pc_mux_sel
+ rst 28 30
+ ICV_30 $T=0 0 0 0 $X=0 $Y=77000
X7 mem_mux_sel<0> dmem_rdata<16> dmem_rdata<15> dmem_rdata<7> 31 33 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<16> imm<15> dmem_addr<16> dmem_addr<15> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30>
+ rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23>
+ rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17>
+ rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10>
+ rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3>
+ rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> rs2_sel<2> rd_sel<1> rs1_sel<1> shift_out<83> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk shift_out<78> shift_out<102> shift_out98> dmem_wdata<16> dmem_wdata<15> shift_out<82> shift_out<77> alu_mux_1_sel
+ imem_addr<10> alu_inv_rs2 alu_mux_2_sel 374 395 shift_out<62> alu_op<0> alu_op<1> shift_dir shift_out<75> shift_out<70> shift_out<85> shift_out<80> shift_out<71> shift_out<42> shift_out<91> shift_out<86> shift_out<57> shift_out<43> shift_out<38>
+ shift_out<123> shift_out<117> shift_out<4> shift_msb shift_out<159> shift_amount<0> shift_out<84> shift_out<81> shift_out<52> shift_amount<1> shift_amount<2> shift_amount<3> shift_out<79> shift_amount<4> cmp_mux_sel 405 384 406 385 386
+ 407 pc_mux_sel rst 32 34
+ ICV_31 $T=0 0 0 0 $X=0 $Y=67600
X8 mem_mux_sel<0> dmem_rdata<20> dmem_rdata<19> dmem_rdata<18> dmem_rdata<17> dmem_rdata<7> dmem_rdata<15> 35 37 39 41 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<20> imm<19> imm<18> imm<17> dmem_addr<20> dmem_addr<19>
+ dmem_addr<18> dmem_addr<17> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26>
+ rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20>
+ rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13>
+ rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6>
+ rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out98> shift_out<92> rs2_sel<2> rd_sel<1> rs1_sel<1> shift_out<87> shift_out<117>
+ shift_out<112> rs2_sel<1> rs2_sel<0> rs1_sel<0> shift_out<107> clk dmem_wdata<20> dmem_wdata<19> dmem_wdata<18> dmem_wdata<17> alu_mux_1_sel imem_addr<10> alu_inv_rs2 alu_mux_2_sel 395 423 shift_out<82> shift_out<72> shift_out<77> alu_op<0>
+ alu_op<1> shift_dir shift_out<95> shift_out<90> shift_out<85> shift_out<80> shift_out<105> shift_out<100> shift_out<91> shift_out<86> shift_out<81> shift_out<52> shift_out<111> shift_out<106> shift_out<101> shift_out<96> shift_out<67> shift_out<122> shift_out<63> shift_out<58>
+ shift_out<53> shift_out<48> shift_out<143> shift_out<138> shift_out<133> shift_out<128> shift_out<24> shift_out<19> shift_out<14> shift_out<9> shift_msb shift_amount<0> shift_amount<1> shift_out<102> shift_amount<2> shift_amount<3> shift_out<104> shift_out<99> shift_out<94> shift_out<89>
+ shift_amount<4> cmp_mux_sel 438 405 439 406 407 440 pc_mux_sel rst 36 38 40 42
+ ICV_36 $T=0 0 0 0 $X=0 $Y=50930
X9 mem_mux_sel<0> dmem_rdata<22> dmem_rdata<21> dmem_rdata<7> dmem_rdata<15> 43 45 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<22> imm<21> dmem_addr<22> dmem_addr<21> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out<107> shift_out<127> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<22> dmem_wdata<21> alu_mux_1_sel imem_addr<22> imem_addr<10> alu_inv_rs2
+ alu_mux_2_sel 449 shift_out<87> shift_out<92> alu_op<0> alu_op<1> shift_dir shift_out<105> shift_out<100> shift_out<115> shift_out<110> shift_out<101> shift_out<96> shift_out<121> shift_out<116> shift_out<132> shift_out<73> shift_out<68> shift_out<153> shift_out<148>
+ shift_out<29> shift_msb shift_amount<0> shift_out<111> shift_out<106> shift_amount<1> shift_out<112> shift_amount<2> shift_amount<3> shift_out<114> shift_out<109> shift_amount<4> cmp_mux_sel 72 438 73 439 440 459 pc_mux_sel
+ rst 44 46
+ ICV_37 $T=0 0 0 0 $X=0 $Y=41600
X10 mem_mux_sel<0> dmem_rdata<24> dmem_rdata<23> dmem_rdata<7> dmem_rdata<15> 47 49 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<24> imm<23> dmem_addr<24> dmem_addr<23> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out<117> shift_out<137> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<24> dmem_wdata<23> alu_mux_1_sel imem_addr<24> imem_addr<23> alu_inv_rs2
+ alu_mux_2_sel 449 469 450 shift_out98> alu_op<0> alu_op<1> shift_dir shift_out<115> shift_out<110> shift_out<125> shift_out<120> shift_out<111> shift_out<106> shift_out<131> shift_out<126> shift_out<142> shift_out<83> shift_out<78> shift_msb
+ shift_out<158> shift_out<44> shift_out<39> shift_amount<0> shift_out<121> shift_out<116> shift_amount<1> shift_out<122> shift_amount<2> shift_out<123> shift_amount<3> shift_out<124> shift_out<119> shift_amount<4> cmp_mux_sel 477 72 74 73 459
+ 478 pc_mux_sel rst 48 50
+ ICV_38 $T=0 0 0 0 $X=0 $Y=32400
X11 mem_mux_sel<0> dmem_rdata<26> dmem_rdata<25> dmem_rdata<7> dmem_rdata<15> 51 53 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<26> imm<25> dmem_addr<26> dmem_addr<25> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out<127> rs2_sel<2> rd_sel<1> rs1_sel<1> rs2_sel<1> rs2_sel<0> rs1_sel<0> shift_out<128> clk dmem_wdata<26> dmem_wdata<25> alu_mux_1_sel imem_addr<26> imem_addr<25> alu_inv_rs2
+ alu_mux_2_sel 487 shift_out<107> shift_out<112> alu_op<0> alu_op<1> shift_dir shift_out<125> shift_out<120> shift_out<135> shift_out<130> shift_out<121> shift_out<116> shift_out<141> shift_out<136> shift_out<152> shift_out<147> shift_out<92> shift_out<87> shift_msb
+ shift_out<54> shift_out<49> shift_amount<0> shift_out<131> shift_out<126> shift_amount<1> shift_out<132> shift_amount<2> shift_out<133> shift_amount<3> shift_out<134> shift_out<129> shift_amount<4> cmp_mux_sel 496 477 497 74 478 498
+ pc_mux_sel rst 52 54
+ ICV_39 $T=0 0 0 0 $X=0 $Y=23150
X12 mem_mux_sel<0> dmem_rdata<28> dmem_rdata<27> dmem_rdata<7> dmem_rdata<15> 55 57 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<28> imm<27> dmem_addr<28> dmem_addr<27> rd_mux_sel<1> rd_mux_sel<2> rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30>
+ rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25> rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24>
+ rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18> rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17>
+ rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12> rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10>
+ rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5> rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4>
+ rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out<137> rs2_sel<2> rd_sel<1> rs1_sel<1> shift_out<138> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk dmem_wdata<28> dmem_wdata<27> alu_mux_1_sel imem_addr<28> imem_addr<27> alu_inv_rs2
+ alu_mux_2_sel 487 507 shift_out<122> shift_out<117> alu_op<0> alu_op<1> shift_dir shift_out<135> shift_out<130> shift_out<145> shift_out<140> shift_out<131> shift_out<126> shift_out<151> shift_out<146> shift_msb shift_out<157> shift_out<102> shift_out98>
+ shift_out<64> shift_out<59> shift_amount<0> shift_out<141> shift_out<136> shift_amount<1> shift_out<142> shift_amount<2> shift_out<143> shift_amount<3> shift_out<144> shift_out<139> shift_amount<4> cmp_mux_sel 515 496 75 497 498 516
+ pc_mux_sel rst 56 58
+ ICV_40 $T=0 0 0 0 $X=0 $Y=13800
X13 mem_mux_sel<0> dmem_rdata<31> dmem_rdata<30> dmem_rdata<29> dmem_rdata<7> dmem_rdata<15> vss! 61 63 mem_mux_sel<1> mem_mux_sel<2> rd_mux_sel<0> imm<31> imm<30> imm<29> dmem_addr<31> dmem_addr<30> dmem_addr<29> rd_mux_sel<1> rd_mux_sel<2>
+ rd_sel<31> rs1_sel<31> rs2_sel<31> rd_sel<30> rs1_sel<30> rs2_sel<30> rd_sel<29> rs1_sel<29> rs2_sel<29> rd_sel<28> rs1_sel<28> rs2_sel<28> rd_sel<27> rs1_sel<27> rs2_sel<27> rd_sel<26> rs1_sel<26> rs2_sel<26> rd_sel<25> rs1_sel<25>
+ rs2_sel<25> rd_sel<24> rs1_sel<24> rs2_sel<24> rd_sel<23> rs1_sel<23> rs2_sel<23> rd_sel<22> rs1_sel<22> rs2_sel<22> rd_sel<21> rs1_sel<21> rs2_sel<21> rd_sel<20> rs1_sel<20> rs2_sel<20> rd_sel<19> rs1_sel<19> rs2_sel<19> rd_sel<18>
+ rs1_sel<18> rs2_sel<18> rd_sel<17> rs1_sel<17> rs2_sel<17> rd_sel<16> rs1_sel<16> rs2_sel<16> rd_sel<15> rs1_sel<15> rs2_sel<15> rd_sel<14> rs1_sel<14> rs2_sel<14> rd_sel<13> rs1_sel<13> rs2_sel<13> rd_sel<12> rs1_sel<12> rs2_sel<12>
+ rd_sel<11> rs1_sel<11> rs2_sel<11> rd_sel<10> rs1_sel<10> rs2_sel<10> rd_sel<9> rs1_sel<9> rs2_sel<9> rd_sel<8> rs1_sel<8> rs2_sel<8> rd_sel<7> rs1_sel<7> rs2_sel<7> rd_sel<6> rs1_sel<6> rs2_sel<6> rd_sel<5> rs1_sel<5>
+ rs2_sel<5> rd_sel<4> rs1_sel<4> rs2_sel<4> rd_sel<3> rs1_sel<3> rs2_sel<3> rd_sel<2> rs1_sel<2> shift_out<148> shift_out<158> rs2_sel<2> rd_sel<1> rs1_sel<1> shift_out<153> rs2_sel<1> rs2_sel<0> rs1_sel<0> clk cmp_a_31
+ dmem_wdata<31> dmem_wdata<30> dmem_wdata<29> alu_mux_1_sel imem_addr<31> imem_addr<30> imem_addr<29> alu_inv_rs2 alu_mux_2_sel shift_out<127> shift_out<132> shift_out<137> alu_op<0> alu_op<1> shift_dir shift_out<150> shift_out<145> shift_out<140> shift_msb shift_out<155>
+ shift_out<146> shift_out<141> shift_out<136> shift_out<156> shift_out<117> shift_out<112> shift_out<107> shift_out<79> shift_out<74> shift_out<69> shift_amount<0> shift_out<151> shift_amount<1> shift_out<157> shift_out<152> shift_out<147> shift_amount<2> shift_amount<3> shift_out<159> shift_out<154>
+ shift_out<149> shift_amount<4> cmp_mux_sel cmp_b_31 60 515 75 516 pc_mux_sel rst 62 64
+ ICV_41 $T=0 0 0 0 $X=0 $Y=0
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
