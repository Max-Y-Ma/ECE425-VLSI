* SPICE NETLIST
***************************************

.SUBCKT bit1 W R A vss! vdd! Z
** N=11 EP=6 IP=0 FDC=14
M0 vss! W 1 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 4 R vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=690 $Y=600 $D=1
M2 5 W A vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=1425 $Y=600 $D=1
M3 vss! 5 8 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=2160 $Y=600 $D=1
M4 6 8 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=2540 $Y=600 $D=1
M5 5 1 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=2985 $Y=600 $D=1
M6 Z R 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=3795 $Y=600 $D=1
M7 vdd! W 1 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M8 4 R vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=690 $Y=1850 $D=0
M9 5 1 A vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=1425 $Y=1850 $D=0
M10 vdd! 5 8 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=2160 $Y=1850 $D=0
M11 6 8 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=2540 $Y=1850 $D=0
M12 5 W 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=2985 $Y=1850 $D=0
M13 Z 4 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=3795 $Y=1850 $D=0
.ENDS
***************************************
