VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  SPACING 0.065 SAMENET ;
  RESISTANCE RPERSQ 0.38 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
  PROPERTY contactResistance 5.69 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.4 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

SITE CoreSite
  CLASS CORE ;
  SIZE 0.005 BY 1.3075 ;
END CoreSite

MACRO aoi21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN aoi21 0 0.1 ;
  SIZE 0.7525 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.085 0.5975 0.15 0.7325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3025 0.5975 0.3675 0.7325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.565 0.49 0.7 0.555 ;
    END
  END C
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6325 0.62 0.6975 1.2425 ;
        RECT 0.4325 0.62 0.6975 0.685 ;
        RECT 0.4325 0.265 0.4975 0.685 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.7525 1.5075 ;
        RECT 0.2425 0.8125 0.3075 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.7525 0.2 ;
        RECT 0.6325 0 0.6975 0.425 ;
        RECT 0.055 0 0.12 0.515 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.4325 0.8125 0.4975 1.2425 ;
      RECT 0.055 0.8125 0.12 1.2425 ;
    LAYER metal2 ;
      RECT 0.43 0.96 0.5 1.095 ;
      RECT 0.0525 0.96 0.1225 1.095 ;
      RECT 0.0525 0.9925 0.5 1.0625 ;
    LAYER via1 ;
      RECT 0.4325 0.995 0.4975 1.06 ;
      RECT 0.055 0.995 0.12 1.06 ;
  END
END aoi21

MACRO buf
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN buf 0 0.1 ;
  SIZE 0.55 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185 0.7925 0.25 0.9275 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.265 0.495 1.2425 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.55 1.5075 ;
        RECT 0.2425 0.9925 0.3075 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.55 0.2 ;
        RECT 0.2425 0 0.3075 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.295 0.5925 0.36 0.7275 ;
      RECT 0.055 0.265 0.12 1.2425 ;
    LAYER metal2 ;
      RECT 0.2925 0.5925 0.3625 0.7275 ;
      RECT 0.0525 0.5925 0.1225 0.7275 ;
      RECT 0.0525 0.625 0.3625 0.695 ;
    LAYER via1 ;
      RECT 0.295 0.6275 0.36 0.6925 ;
      RECT 0.055 0.6275 0.12 0.6925 ;
  END
END buf

MACRO dff
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN dff 0 0.1 ;
  SIZE 4.3425 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.04 0.6 0.175 0.665 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7 0.5975 0.835 0.6625 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.46 0.265 3.525 1.2425 ;
    END
  END Q
  PIN Qb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.095 0.745 3.725 0.815 ;
      LAYER metal1 ;
        RECT 3.59 0.7475 3.725 0.8125 ;
        RECT 3.13 0.55 3.395 0.615 ;
        RECT 3.095 0.7475 3.23 0.8125 ;
        RECT 3.13 0.265 3.195 1.2425 ;
      LAYER via1 ;
        RECT 3.13 0.7475 3.195 0.8125 ;
        RECT 3.625 0.7475 3.69 0.8125 ;
    END
  END Qb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 4.3425 1.5075 ;
        RECT 3.605 0.9925 3.67 1.5075 ;
        RECT 3.275 0.9925 3.34 1.5075 ;
        RECT 2.945 0.9925 3.01 1.5075 ;
        RECT 1.8075 0.9925 1.8725 1.5075 ;
        RECT 1.4775 0.9925 1.5425 1.5075 ;
        RECT 0.715 0.9925 0.78 1.5075 ;
        RECT 0.385 0.9925 0.45 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 4.3425 0.2 ;
        RECT 3.605 0 3.67 0.425 ;
        RECT 3.275 0 3.34 0.425 ;
        RECT 2.945 0 3.01 0.425 ;
        RECT 1.8075 0 1.8725 0.425 ;
        RECT 1.4775 0 1.5425 0.425 ;
        RECT 0.715 0 0.78 0.425 ;
        RECT 0.385 0 0.45 0.425 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 4.2225 0.265 4.2875 1.2425 ;
      RECT 4.1875 0.6075 4.3225 0.6725 ;
      RECT 2.7975 0.265 2.8625 1.2425 ;
      RECT 2.6925 0.6075 2.8625 0.6725 ;
      RECT 2.7975 0.55 3.065 0.615 ;
      RECT 2.4675 0.265 2.5325 1.2425 ;
      RECT 2.455 0.7475 2.59 0.8125 ;
      RECT 2.3225 0.265 2.3875 1.2425 ;
      RECT 2.2175 0.6075 2.3875 0.6725 ;
      RECT 1.6625 0.265 1.7275 1.2425 ;
      RECT 1.6275 0.7475 1.7625 0.8125 ;
      RECT 1.6625 0.5275 1.9275 0.5925 ;
      RECT 1.3325 0.265 1.3975 1.2425 ;
      RECT 1.2975 0.6075 1.5975 0.6725 ;
      RECT 0.24 0.265 0.305 1.2425 ;
      RECT 0.24 0.5275 0.505 0.5925 ;
      RECT 4.0225 0.465 4.1575 0.53 ;
      RECT 3.92 0.8875 4.055 0.9525 ;
      RECT 3.79 0.265 3.855 1.2425 ;
      RECT 2.5975 0.465 2.7325 0.53 ;
      RECT 2.5975 0.8875 2.7325 0.9525 ;
      RECT 2.1225 0.465 2.2575 0.53 ;
      RECT 2.1225 0.8875 2.2575 0.9525 ;
      RECT 1.9925 0.265 2.0575 1.2425 ;
      RECT 1.1325 0.4675 1.2675 0.5325 ;
      RECT 1.03 0.8875 1.165 0.9525 ;
      RECT 0.9 0.265 0.965 1.2425 ;
      RECT 0.57 0.265 0.635 1.2425 ;
    LAYER metal2 ;
      RECT 0.5675 0.43 0.6375 0.565 ;
      RECT 1.1325 0.4625 1.2675 0.535 ;
      RECT 0.5675 0.4625 4.1575 0.5325 ;
      RECT 0.2375 0.855 0.3075 0.99 ;
      RECT 0.2375 0.885 4.055 0.955 ;
      RECT 2.6925 0.605 4.3225 0.675 ;
      RECT 1.6275 0.745 2.59 0.815 ;
      RECT 1.2975 0.605 2.3525 0.675 ;
    LAYER via1 ;
      RECT 4.2225 0.6075 4.2875 0.6725 ;
      RECT 4.0575 0.465 4.1225 0.53 ;
      RECT 3.955 0.8875 4.02 0.9525 ;
      RECT 2.7275 0.6075 2.7925 0.6725 ;
      RECT 2.6325 0.465 2.6975 0.53 ;
      RECT 2.6325 0.8875 2.6975 0.9525 ;
      RECT 2.49 0.7475 2.555 0.8125 ;
      RECT 2.2525 0.6075 2.3175 0.6725 ;
      RECT 2.1575 0.465 2.2225 0.53 ;
      RECT 2.1575 0.8875 2.2225 0.9525 ;
      RECT 1.6625 0.7475 1.7275 0.8125 ;
      RECT 1.3325 0.6075 1.3975 0.6725 ;
      RECT 1.1675 0.4675 1.2325 0.5325 ;
      RECT 1.065 0.8875 1.13 0.9525 ;
      RECT 0.57 0.465 0.635 0.53 ;
      RECT 0.24 0.89 0.305 0.955 ;
  END
END dff

MACRO dlatch
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN dlatch 0 0.1 ;
  SIZE 2.4425 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7 0.655 0.835 0.72 ;
    END
  END D
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.04 0.655 0.175 0.72 ;
    END
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.56 0.7225 1.825 0.7875 ;
        RECT 1.56 0.265 1.625 1.2425 ;
    END
  END Q
  PIN Qb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.89 0.265 1.955 1.2425 ;
    END
  END Qb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 2.4425 1.5075 ;
        RECT 1.705 0.9925 1.77 1.5075 ;
        RECT 1.375 0.9925 1.44 1.5075 ;
        RECT 0.715 0.9925 0.78 1.5075 ;
        RECT 0.385 0.9925 0.45 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 2.4425 0.2 ;
        RECT 1.705 0 1.77 0.425 ;
        RECT 1.375 0 1.44 0.425 ;
        RECT 0.715 0 0.78 0.425 ;
        RECT 0.385 0 0.45 0.425 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 1.23 0.265 1.295 1.2425 ;
      RECT 1.23 0.6075 1.495 0.6725 ;
      RECT 0.24 0.265 0.305 1.2425 ;
      RECT 0.24 0.655 0.505 0.72 ;
      RECT 2.3225 0.265 2.3875 1.2425 ;
      RECT 2.1225 0.465 2.2575 0.53 ;
      RECT 2.02 0.8875 2.155 0.9525 ;
      RECT 1.03 0.465 1.165 0.53 ;
      RECT 1.03 0.8875 1.165 0.9525 ;
      RECT 0.9 0.265 0.965 1.2425 ;
      RECT 0.57 0.265 0.635 1.2425 ;
    LAYER metal2 ;
      RECT 2.32 0.5725 2.39 0.7075 ;
      RECT 1.2975 0.605 2.39 0.675 ;
      RECT 0.5675 0.43 0.6375 0.565 ;
      RECT 0.5675 0.4625 2.2575 0.5325 ;
      RECT 0.2375 0.855 0.3075 0.99 ;
      RECT 0.2375 0.885 2.155 0.955 ;
    LAYER via1 ;
      RECT 2.3225 0.6075 2.3875 0.6725 ;
      RECT 2.1575 0.465 2.2225 0.53 ;
      RECT 2.055 0.8875 2.12 0.9525 ;
      RECT 1.3325 0.6075 1.3975 0.6725 ;
      RECT 1.065 0.465 1.13 0.53 ;
      RECT 1.065 0.8875 1.13 0.9525 ;
      RECT 0.57 0.465 0.635 0.53 ;
      RECT 0.24 0.89 0.305 0.955 ;
  END
END dlatch

MACRO inv
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN inv 0 0.1 ;
  SIZE 0.36 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.04 0.655 0.175 0.72 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.24 0.265 0.305 1.2425 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.36 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.36 0.2 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
END inv

MACRO mux2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN mux2 0 0.1 ;
  SIZE 1.625 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615 0.5825 0.68 0.7175 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.91 0.5525 1.045 0.6175 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.0825 0.5775 1.245 0.6475 ;
        RECT 0.0825 0.545 0.1525 0.68 ;
      LAYER metal1 ;
        RECT 1.11 0.58 1.245 0.645 ;
        RECT 0.085 0.545 0.15 0.68 ;
      LAYER via1 ;
        RECT 0.085 0.58 0.15 0.645 ;
        RECT 1.145 0.58 1.21 0.645 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.505 0.265 1.57 1.2425 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 1.625 1.5075 ;
        RECT 1.32 0.9925 1.385 1.5075 ;
        RECT 0.5725 0.8125 0.6375 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.625 0.2 ;
        RECT 1.32 0 1.385 0.425 ;
        RECT 1.175 0 1.24 0.515 ;
        RECT 0.385 0 0.45 0.515 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.9875 0.6825 1.0525 1.2425 ;
      RECT 0.9525 0.72 1.0875 0.785 ;
      RECT 0.78 0.6825 1.0525 0.7475 ;
      RECT 0.78 0.265 0.845 0.7475 ;
      RECT 0.24 0.265 0.305 1.2425 ;
      RECT 0.24 0.65 0.505 0.715 ;
      RECT 1.305 0.72 1.44 0.785 ;
      RECT 1.175 0.8125 1.24 1.2425 ;
      RECT 0.78 0.8125 0.845 1.2425 ;
      RECT 0.385 0.8125 0.45 1.2425 ;
    LAYER metal2 ;
      RECT 1.1725 0.9925 1.2425 1.1275 ;
      RECT 0.7775 0.9925 0.8475 1.1275 ;
      RECT 0.3825 0.9925 0.4525 1.1275 ;
      RECT 0.3825 1.025 1.2425 1.095 ;
      RECT 0.9525 0.7175 1.44 0.7875 ;
    LAYER via1 ;
      RECT 1.34 0.72 1.405 0.785 ;
      RECT 1.175 1.0275 1.24 1.0925 ;
      RECT 0.9875 0.72 1.0525 0.785 ;
      RECT 0.78 1.0275 0.845 1.0925 ;
      RECT 0.385 1.0275 0.45 1.0925 ;
  END
END mux2

MACRO nand2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nand2 0 0.1 ;
  SIZE 0.55 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.04 0.575 0.175 0.64 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.41 0.71 0.475 0.845 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2425 0.575 0.495 0.64 ;
        RECT 0.43 0.265 0.495 0.64 ;
        RECT 0.2425 0.575 0.3075 1.2425 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.55 1.5075 ;
        RECT 0.43 0.9925 0.495 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.55 0.2 ;
        RECT 0.055 0 0.12 0.515 ;
    END
  END vss!
END nand2

MACRO nor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nor2 0 0.1 ;
  SIZE 0.55 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.04 0.575 0.175 0.64 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4 0.49 0.465 0.625 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.69 0.495 1.2425 ;
        RECT 0.2425 0.69 0.495 0.755 ;
        RECT 0.2425 0.265 0.3075 0.755 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.55 1.5075 ;
        RECT 0.055 0.8125 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.55 0.2 ;
        RECT 0.43 0 0.495 0.425 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
END nor2

MACRO oai21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN oai21 0 0.1 ;
  SIZE 0.76 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0425 0.6825 0.1775 0.7475 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3725 0.585 0.5075 0.65 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5725 0.715 0.7075 0.78 ;
    END
  END C
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.715 0.495 1.2425 ;
        RECT 0.2425 0.715 0.495 0.78 ;
        RECT 0.2425 0.265 0.3075 0.78 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.76 1.5075 ;
        RECT 0.64 0.9925 0.705 1.5075 ;
        RECT 0.055 0.8125 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.76 0.2 ;
        RECT 0.64 0 0.705 0.515 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.43 0.265 0.495 0.515 ;
      RECT 0.055 0.265 0.12 0.515 ;
    LAYER metal2 ;
      RECT 0.4275 0.3225 0.4975 0.4575 ;
      RECT 0.0525 0.3225 0.1225 0.4575 ;
      RECT 0.0525 0.355 0.4975 0.425 ;
    LAYER via1 ;
      RECT 0.43 0.3575 0.495 0.4225 ;
      RECT 0.055 0.3575 0.12 0.4225 ;
  END
END oai21

MACRO or2
  CLASS CORE ;
  ORIGIN 0 -0.1025 ;
  FOREIGN or2 0 0.1025 ;
  SIZE 0.76 BY 1.305 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.035 0.5275 0.17 0.5925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3725 0.49 0.5075 0.555 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.64 0.265 0.705 1.2425 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 0.76 1.5075 ;
        RECT 0.43 0.8125 0.495 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.76 0.2 ;
        RECT 0.43 0 0.495 0.425 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.055 0.68 0.12 1.2425 ;
      RECT 0.055 0.68 0.575 0.745 ;
      RECT 0.2425 0.265 0.3075 0.745 ;
  END
END or2

MACRO xnor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xnor2 0 0.1 ;
  SIZE 1.28 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.04 0.5775 0.6975 0.6475 ;
      LAYER metal1 ;
        RECT 0.5625 0.58 0.6975 0.645 ;
        RECT 0.04 0.58 0.175 0.645 ;
      LAYER via1 ;
        RECT 0.075 0.58 0.14 0.645 ;
        RECT 0.5975 0.58 0.6625 0.645 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.8925 0.5825 1.0275 0.6525 ;
        RECT 0.4075 0.75 0.995 0.82 ;
        RECT 0.925 0.5825 0.995 0.82 ;
        RECT 0.4075 0.7175 0.4775 0.8525 ;
      LAYER metal1 ;
        RECT 0.8925 0.585 1.0275 0.65 ;
        RECT 0.41 0.7175 0.475 0.8525 ;
      LAYER via1 ;
        RECT 0.41 0.7525 0.475 0.8175 ;
        RECT 0.9275 0.585 0.9925 0.65 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.95 0.715 1.015 1.2425 ;
        RECT 0.7625 0.715 1.015 0.78 ;
        RECT 0.7625 0.265 0.8275 0.78 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 1.28 1.5075 ;
        RECT 1.16 0.9925 1.225 1.5075 ;
        RECT 0.575 0.8125 0.64 1.5075 ;
        RECT 0.43 0.9925 0.495 1.5075 ;
        RECT 0.055 0.9925 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.28 0.2 ;
        RECT 1.16 0 1.225 0.515 ;
        RECT 0.055 0 0.12 0.515 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.2425 0.575 0.3075 1.2425 ;
      RECT 0.2425 0.575 0.495 0.64 ;
      RECT 0.43 0.265 0.495 0.64 ;
      RECT 1.0925 0.765 1.2275 0.83 ;
      RECT 0.95 0.265 1.015 0.515 ;
      RECT 0.575 0.265 0.64 0.515 ;
    LAYER metal2 ;
      RECT 0.24 0.89 0.31 1.025 ;
      RECT 0.24 0.9225 1.1975 0.9925 ;
      RECT 1.1275 0.7625 1.1975 0.9925 ;
      RECT 1.0925 0.7625 1.2275 0.8325 ;
      RECT 0.9475 0.3225 1.0175 0.4575 ;
      RECT 0.5725 0.3225 0.6425 0.4575 ;
      RECT 0.5725 0.355 1.0175 0.425 ;
    LAYER via1 ;
      RECT 1.1275 0.765 1.1925 0.83 ;
      RECT 0.95 0.3575 1.015 0.4225 ;
      RECT 0.575 0.3575 0.64 0.4225 ;
      RECT 0.2425 0.925 0.3075 0.99 ;
  END
END xnor2

MACRO xor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xor2 0 0.1 ;
  SIZE 1.275 BY 1.3075 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.0725 0.745 0.6775 0.815 ;
        RECT 0.6075 0.5975 0.6775 0.815 ;
        RECT 0.04 0.5725 0.175 0.6425 ;
        RECT 0.0725 0.5725 0.1425 0.815 ;
      LAYER metal1 ;
        RECT 0.61 0.5975 0.675 0.7325 ;
        RECT 0.04 0.575 0.175 0.64 ;
      LAYER via1 ;
        RECT 0.075 0.575 0.14 0.64 ;
        RECT 0.61 0.6325 0.675 0.6975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.8225 0.435 0.8925 0.7325 ;
        RECT 0.3975 0.435 0.8925 0.505 ;
        RECT 0.3975 0.435 0.4675 0.625 ;
      LAYER metal1 ;
        RECT 0.825 0.5975 0.89 0.7325 ;
        RECT 0.4 0.49 0.465 0.625 ;
      LAYER via1 ;
        RECT 0.4 0.525 0.465 0.59 ;
        RECT 0.825 0.6325 0.89 0.6975 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.155 0.62 1.22 1.2425 ;
        RECT 0.955 0.62 1.22 0.685 ;
        RECT 0.955 0.265 1.02 0.685 ;
    END
  END Z
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.3075 1.275 1.5075 ;
        RECT 0.765 0.8125 0.83 1.5075 ;
        RECT 0.055 0.8125 0.12 1.5075 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.275 0.2 ;
        RECT 1.155 0 1.22 0.425 ;
        RECT 0.5775 0 0.6425 0.515 ;
        RECT 0.43 0 0.495 0.425 ;
        RECT 0.055 0 0.12 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.43 0.69 0.495 1.2425 ;
      RECT 0.2425 0.69 0.495 0.755 ;
      RECT 0.2425 0.265 0.3075 0.755 ;
      RECT 1.0875 0.49 1.2225 0.555 ;
      RECT 0.955 0.8125 1.02 1.2425 ;
      RECT 0.5775 0.8125 0.6425 1.2425 ;
    LAYER metal2 ;
      RECT 1.0875 0.4875 1.2225 0.5575 ;
      RECT 0.24 0.295 0.31 0.5425 ;
      RECT 1.12 0.295 1.19 0.5575 ;
      RECT 0.24 0.295 1.19 0.365 ;
      RECT 0.9525 0.96 1.0225 1.095 ;
      RECT 0.575 0.96 0.645 1.095 ;
      RECT 0.575 0.9925 1.0225 1.0625 ;
    LAYER via1 ;
      RECT 1.1225 0.49 1.1875 0.555 ;
      RECT 0.955 0.995 1.02 1.06 ;
      RECT 0.5775 0.995 0.6425 1.06 ;
      RECT 0.2425 0.4425 0.3075 0.5075 ;
  END
END xor2

MACRO regfile
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN regfile 0 0 ;
  SIZE 88.91 BY 1.405 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.1725 0.975 87.24 1.045 ;
        RECT 87.17 0.69 87.24 1.045 ;
        RECT 85.1725 0.69 85.2425 1.045 ;
      LAYER metal1 ;
        RECT 87.1725 0.69 87.2475 0.825 ;
        RECT 85.175 0.69 85.25 0.825 ;
      LAYER via1 ;
        RECT 85.175 0.725 85.24 0.79 ;
        RECT 87.1725 0.725 87.2375 0.79 ;
    END
  END clk
  PIN rd_mux_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.575 0.2625 81.71 0.3325 ;
        RECT 81.6075 0.115 81.6775 0.3325 ;
        RECT 0.6075 0.115 81.6775 0.185 ;
        RECT 78.875 0.2625 79.01 0.3325 ;
        RECT 78.9075 0.115 78.9775 0.3325 ;
        RECT 76.175 0.2625 76.31 0.3325 ;
        RECT 76.2075 0.115 76.2775 0.3325 ;
        RECT 73.475 0.2625 73.61 0.3325 ;
        RECT 73.5075 0.115 73.5775 0.3325 ;
        RECT 70.775 0.2625 70.91 0.3325 ;
        RECT 70.8075 0.115 70.8775 0.3325 ;
        RECT 68.075 0.2625 68.21 0.3325 ;
        RECT 68.1075 0.115 68.1775 0.3325 ;
        RECT 65.375 0.2625 65.51 0.3325 ;
        RECT 65.4075 0.115 65.4775 0.3325 ;
        RECT 62.675 0.2625 62.81 0.3325 ;
        RECT 62.7075 0.115 62.7775 0.3325 ;
        RECT 59.975 0.2625 60.11 0.3325 ;
        RECT 60.0075 0.115 60.0775 0.3325 ;
        RECT 57.275 0.2625 57.41 0.3325 ;
        RECT 57.3075 0.115 57.3775 0.3325 ;
        RECT 54.575 0.2625 54.71 0.3325 ;
        RECT 54.6075 0.115 54.6775 0.3325 ;
        RECT 51.875 0.2625 52.01 0.3325 ;
        RECT 51.9075 0.115 51.9775 0.3325 ;
        RECT 49.175 0.2625 49.31 0.3325 ;
        RECT 49.2075 0.115 49.2775 0.3325 ;
        RECT 46.475 0.2625 46.61 0.3325 ;
        RECT 46.5075 0.115 46.5775 0.3325 ;
        RECT 43.775 0.2625 43.91 0.3325 ;
        RECT 43.8075 0.115 43.8775 0.3325 ;
        RECT 41.075 0.2625 41.21 0.3325 ;
        RECT 41.1075 0.115 41.1775 0.3325 ;
        RECT 38.375 0.2625 38.51 0.3325 ;
        RECT 38.4075 0.115 38.4775 0.3325 ;
        RECT 35.675 0.2625 35.81 0.3325 ;
        RECT 35.7075 0.115 35.7775 0.3325 ;
        RECT 32.975 0.2625 33.11 0.3325 ;
        RECT 33.0075 0.115 33.0775 0.3325 ;
        RECT 30.275 0.2625 30.41 0.3325 ;
        RECT 30.3075 0.115 30.3775 0.3325 ;
        RECT 27.575 0.2625 27.71 0.3325 ;
        RECT 27.6075 0.115 27.6775 0.3325 ;
        RECT 24.875 0.2625 25.01 0.3325 ;
        RECT 24.9075 0.115 24.9775 0.3325 ;
        RECT 22.175 0.2625 22.31 0.3325 ;
        RECT 22.2075 0.115 22.2775 0.3325 ;
        RECT 19.475 0.2625 19.61 0.3325 ;
        RECT 19.5075 0.115 19.5775 0.3325 ;
        RECT 16.775 0.2625 16.91 0.3325 ;
        RECT 16.8075 0.115 16.8775 0.3325 ;
        RECT 14.075 0.2625 14.21 0.3325 ;
        RECT 14.1075 0.115 14.1775 0.3325 ;
        RECT 11.375 0.2625 11.51 0.3325 ;
        RECT 11.4075 0.115 11.4775 0.3325 ;
        RECT 8.675 0.2625 8.81 0.3325 ;
        RECT 8.7075 0.115 8.7775 0.3325 ;
        RECT 5.975 0.2625 6.11 0.3325 ;
        RECT 6.0075 0.115 6.0775 0.3325 ;
        RECT 3.275 0.2625 3.41 0.3325 ;
        RECT 3.3075 0.115 3.3775 0.3325 ;
        RECT 0.575 0.2625 0.71 0.3325 ;
        RECT 0.6075 0.115 0.6775 0.3325 ;
      LAYER metal1 ;
        RECT 81.575 0.265 81.71 0.33 ;
        RECT 81.575 0.265 81.64 1.14 ;
        RECT 78.875 0.265 79.01 0.33 ;
        RECT 78.875 0.265 78.94 1.14 ;
        RECT 76.175 0.265 76.31 0.33 ;
        RECT 76.175 0.265 76.24 1.14 ;
        RECT 73.475 0.265 73.61 0.33 ;
        RECT 73.475 0.265 73.54 1.14 ;
        RECT 70.775 0.265 70.91 0.33 ;
        RECT 70.775 0.265 70.84 1.14 ;
        RECT 68.075 0.265 68.21 0.33 ;
        RECT 68.075 0.265 68.14 1.14 ;
        RECT 65.375 0.265 65.51 0.33 ;
        RECT 65.375 0.265 65.44 1.14 ;
        RECT 62.675 0.265 62.81 0.33 ;
        RECT 62.675 0.265 62.74 1.14 ;
        RECT 59.975 0.265 60.11 0.33 ;
        RECT 59.975 0.265 60.04 1.14 ;
        RECT 57.275 0.265 57.41 0.33 ;
        RECT 57.275 0.265 57.34 1.14 ;
        RECT 54.575 0.265 54.71 0.33 ;
        RECT 54.575 0.265 54.64 1.14 ;
        RECT 51.875 0.265 52.01 0.33 ;
        RECT 51.875 0.265 51.94 1.14 ;
        RECT 49.175 0.265 49.31 0.33 ;
        RECT 49.175 0.265 49.24 1.14 ;
        RECT 46.475 0.265 46.61 0.33 ;
        RECT 46.475 0.265 46.54 1.14 ;
        RECT 43.775 0.265 43.91 0.33 ;
        RECT 43.775 0.265 43.84 1.14 ;
        RECT 41.075 0.265 41.21 0.33 ;
        RECT 41.075 0.265 41.14 1.14 ;
        RECT 38.375 0.265 38.51 0.33 ;
        RECT 38.375 0.265 38.44 1.14 ;
        RECT 35.675 0.265 35.81 0.33 ;
        RECT 35.675 0.265 35.74 1.14 ;
        RECT 32.975 0.265 33.11 0.33 ;
        RECT 32.975 0.265 33.04 1.14 ;
        RECT 30.275 0.265 30.41 0.33 ;
        RECT 30.275 0.265 30.34 1.14 ;
        RECT 27.575 0.265 27.71 0.33 ;
        RECT 27.575 0.265 27.64 1.14 ;
        RECT 24.875 0.265 25.01 0.33 ;
        RECT 24.875 0.265 24.94 1.14 ;
        RECT 22.175 0.265 22.31 0.33 ;
        RECT 22.175 0.265 22.24 1.14 ;
        RECT 19.475 0.265 19.61 0.33 ;
        RECT 19.475 0.265 19.54 1.14 ;
        RECT 16.775 0.265 16.91 0.33 ;
        RECT 16.775 0.265 16.84 1.14 ;
        RECT 14.075 0.265 14.21 0.33 ;
        RECT 14.075 0.265 14.14 1.14 ;
        RECT 11.375 0.265 11.51 0.33 ;
        RECT 11.375 0.265 11.44 1.14 ;
        RECT 8.675 0.265 8.81 0.33 ;
        RECT 8.675 0.265 8.74 1.14 ;
        RECT 5.975 0.265 6.11 0.33 ;
        RECT 5.975 0.265 6.04 1.14 ;
        RECT 3.275 0.265 3.41 0.33 ;
        RECT 3.275 0.265 3.34 1.14 ;
        RECT 0.575 0.265 0.71 0.33 ;
        RECT 0.575 0.265 0.64 1.14 ;
      LAYER via1 ;
        RECT 0.61 0.265 0.675 0.33 ;
        RECT 3.31 0.265 3.375 0.33 ;
        RECT 6.01 0.265 6.075 0.33 ;
        RECT 8.71 0.265 8.775 0.33 ;
        RECT 11.41 0.265 11.475 0.33 ;
        RECT 14.11 0.265 14.175 0.33 ;
        RECT 16.81 0.265 16.875 0.33 ;
        RECT 19.51 0.265 19.575 0.33 ;
        RECT 22.21 0.265 22.275 0.33 ;
        RECT 24.91 0.265 24.975 0.33 ;
        RECT 27.61 0.265 27.675 0.33 ;
        RECT 30.31 0.265 30.375 0.33 ;
        RECT 33.01 0.265 33.075 0.33 ;
        RECT 35.71 0.265 35.775 0.33 ;
        RECT 38.41 0.265 38.475 0.33 ;
        RECT 41.11 0.265 41.175 0.33 ;
        RECT 43.81 0.265 43.875 0.33 ;
        RECT 46.51 0.265 46.575 0.33 ;
        RECT 49.21 0.265 49.275 0.33 ;
        RECT 51.91 0.265 51.975 0.33 ;
        RECT 54.61 0.265 54.675 0.33 ;
        RECT 57.31 0.265 57.375 0.33 ;
        RECT 60.01 0.265 60.075 0.33 ;
        RECT 62.71 0.265 62.775 0.33 ;
        RECT 65.41 0.265 65.475 0.33 ;
        RECT 68.11 0.265 68.175 0.33 ;
        RECT 70.81 0.265 70.875 0.33 ;
        RECT 73.51 0.265 73.575 0.33 ;
        RECT 76.21 0.265 76.275 0.33 ;
        RECT 78.91 0.265 78.975 0.33 ;
        RECT 81.61 0.265 81.675 0.33 ;
    END
  END rd_mux_out
  PIN rd_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 56.885 0.69 57.025 0.76 ;
      LAYER metal2 ;
        RECT 58.1825 0.77 58.2525 0.905 ;
        RECT 58.01 0.77 58.2525 0.84 ;
        RECT 58.01 0.55 58.08 0.84 ;
        RECT 57.25 0.55 58.08 0.62 ;
        RECT 57.4025 0.55 57.4725 0.7 ;
        RECT 56.885 0.69 57.32 0.76 ;
        RECT 57.25 0.55 57.32 0.76 ;
      LAYER metal1 ;
        RECT 58.185 0.77 58.25 0.905 ;
        RECT 57.405 0.565 57.47 0.7 ;
        RECT 56.885 0.6925 57.02 0.7575 ;
        RECT 56.885 0.69 56.95 0.825 ;
      LAYER via2 ;
        RECT 56.92 0.69 56.99 0.76 ;
      LAYER via1 ;
        RECT 56.92 0.6925 56.985 0.7575 ;
        RECT 57.405 0.6 57.47 0.665 ;
        RECT 58.185 0.805 58.25 0.87 ;
    END
  END rd_sel[10]
  PIN rd_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 54.185 0.69 54.325 0.76 ;
      LAYER metal2 ;
        RECT 55.4825 0.77 55.5525 0.905 ;
        RECT 55.31 0.77 55.5525 0.84 ;
        RECT 55.31 0.55 55.38 0.84 ;
        RECT 54.55 0.55 55.38 0.62 ;
        RECT 54.7025 0.55 54.7725 0.7 ;
        RECT 54.185 0.69 54.62 0.76 ;
        RECT 54.55 0.55 54.62 0.76 ;
      LAYER metal1 ;
        RECT 55.485 0.77 55.55 0.905 ;
        RECT 54.705 0.565 54.77 0.7 ;
        RECT 54.185 0.6925 54.32 0.7575 ;
        RECT 54.185 0.69 54.25 0.825 ;
      LAYER via2 ;
        RECT 54.22 0.69 54.29 0.76 ;
      LAYER via1 ;
        RECT 54.22 0.6925 54.285 0.7575 ;
        RECT 54.705 0.6 54.77 0.665 ;
        RECT 55.485 0.805 55.55 0.87 ;
    END
  END rd_sel[11]
  PIN rd_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 51.485 0.69 51.625 0.76 ;
      LAYER metal2 ;
        RECT 52.7825 0.77 52.8525 0.905 ;
        RECT 52.61 0.77 52.8525 0.84 ;
        RECT 52.61 0.55 52.68 0.84 ;
        RECT 51.85 0.55 52.68 0.62 ;
        RECT 52.0025 0.55 52.0725 0.7 ;
        RECT 51.485 0.69 51.92 0.76 ;
        RECT 51.85 0.55 51.92 0.76 ;
      LAYER metal1 ;
        RECT 52.785 0.77 52.85 0.905 ;
        RECT 52.005 0.565 52.07 0.7 ;
        RECT 51.485 0.6925 51.62 0.7575 ;
        RECT 51.485 0.69 51.55 0.825 ;
      LAYER via2 ;
        RECT 51.52 0.69 51.59 0.76 ;
      LAYER via1 ;
        RECT 51.52 0.6925 51.585 0.7575 ;
        RECT 52.005 0.6 52.07 0.665 ;
        RECT 52.785 0.805 52.85 0.87 ;
    END
  END rd_sel[12]
  PIN rd_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 48.785 0.69 48.925 0.76 ;
      LAYER metal2 ;
        RECT 50.0825 0.77 50.1525 0.905 ;
        RECT 49.91 0.77 50.1525 0.84 ;
        RECT 49.91 0.55 49.98 0.84 ;
        RECT 49.15 0.55 49.98 0.62 ;
        RECT 49.3025 0.55 49.3725 0.7 ;
        RECT 48.785 0.69 49.22 0.76 ;
        RECT 49.15 0.55 49.22 0.76 ;
      LAYER metal1 ;
        RECT 50.085 0.77 50.15 0.905 ;
        RECT 49.305 0.565 49.37 0.7 ;
        RECT 48.785 0.6925 48.92 0.7575 ;
        RECT 48.785 0.69 48.85 0.825 ;
      LAYER via2 ;
        RECT 48.82 0.69 48.89 0.76 ;
      LAYER via1 ;
        RECT 48.82 0.6925 48.885 0.7575 ;
        RECT 49.305 0.6 49.37 0.665 ;
        RECT 50.085 0.805 50.15 0.87 ;
    END
  END rd_sel[13]
  PIN rd_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.085 0.69 46.225 0.76 ;
      LAYER metal2 ;
        RECT 47.3825 0.77 47.4525 0.905 ;
        RECT 47.21 0.77 47.4525 0.84 ;
        RECT 47.21 0.55 47.28 0.84 ;
        RECT 46.45 0.55 47.28 0.62 ;
        RECT 46.6025 0.55 46.6725 0.7 ;
        RECT 46.085 0.69 46.52 0.76 ;
        RECT 46.45 0.55 46.52 0.76 ;
      LAYER metal1 ;
        RECT 47.385 0.77 47.45 0.905 ;
        RECT 46.605 0.565 46.67 0.7 ;
        RECT 46.085 0.6925 46.22 0.7575 ;
        RECT 46.085 0.69 46.15 0.825 ;
      LAYER via2 ;
        RECT 46.12 0.69 46.19 0.76 ;
      LAYER via1 ;
        RECT 46.12 0.6925 46.185 0.7575 ;
        RECT 46.605 0.6 46.67 0.665 ;
        RECT 47.385 0.805 47.45 0.87 ;
    END
  END rd_sel[14]
  PIN rd_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 43.385 0.69 43.525 0.76 ;
      LAYER metal2 ;
        RECT 44.6825 0.77 44.7525 0.905 ;
        RECT 44.51 0.77 44.7525 0.84 ;
        RECT 44.51 0.55 44.58 0.84 ;
        RECT 43.75 0.55 44.58 0.62 ;
        RECT 43.9025 0.55 43.9725 0.7 ;
        RECT 43.385 0.69 43.82 0.76 ;
        RECT 43.75 0.55 43.82 0.76 ;
      LAYER metal1 ;
        RECT 44.685 0.77 44.75 0.905 ;
        RECT 43.905 0.565 43.97 0.7 ;
        RECT 43.385 0.6925 43.52 0.7575 ;
        RECT 43.385 0.69 43.45 0.825 ;
      LAYER via2 ;
        RECT 43.42 0.69 43.49 0.76 ;
      LAYER via1 ;
        RECT 43.42 0.6925 43.485 0.7575 ;
        RECT 43.905 0.6 43.97 0.665 ;
        RECT 44.685 0.805 44.75 0.87 ;
    END
  END rd_sel[15]
  PIN rd_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 40.685 0.69 40.825 0.76 ;
      LAYER metal2 ;
        RECT 41.9825 0.77 42.0525 0.905 ;
        RECT 41.81 0.77 42.0525 0.84 ;
        RECT 41.81 0.55 41.88 0.84 ;
        RECT 41.05 0.55 41.88 0.62 ;
        RECT 41.2025 0.55 41.2725 0.7 ;
        RECT 40.685 0.69 41.12 0.76 ;
        RECT 41.05 0.55 41.12 0.76 ;
      LAYER metal1 ;
        RECT 41.985 0.77 42.05 0.905 ;
        RECT 41.205 0.565 41.27 0.7 ;
        RECT 40.685 0.6925 40.82 0.7575 ;
        RECT 40.685 0.69 40.75 0.825 ;
      LAYER via2 ;
        RECT 40.72 0.69 40.79 0.76 ;
      LAYER via1 ;
        RECT 40.72 0.6925 40.785 0.7575 ;
        RECT 41.205 0.6 41.27 0.665 ;
        RECT 41.985 0.805 42.05 0.87 ;
    END
  END rd_sel[16]
  PIN rd_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 37.985 0.69 38.125 0.76 ;
      LAYER metal2 ;
        RECT 39.2825 0.77 39.3525 0.905 ;
        RECT 39.11 0.77 39.3525 0.84 ;
        RECT 39.11 0.55 39.18 0.84 ;
        RECT 38.35 0.55 39.18 0.62 ;
        RECT 38.5025 0.55 38.5725 0.7 ;
        RECT 37.985 0.69 38.42 0.76 ;
        RECT 38.35 0.55 38.42 0.76 ;
      LAYER metal1 ;
        RECT 39.285 0.77 39.35 0.905 ;
        RECT 38.505 0.565 38.57 0.7 ;
        RECT 37.985 0.6925 38.12 0.7575 ;
        RECT 37.985 0.69 38.05 0.825 ;
      LAYER via2 ;
        RECT 38.02 0.69 38.09 0.76 ;
      LAYER via1 ;
        RECT 38.02 0.6925 38.085 0.7575 ;
        RECT 38.505 0.6 38.57 0.665 ;
        RECT 39.285 0.805 39.35 0.87 ;
    END
  END rd_sel[17]
  PIN rd_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 35.285 0.69 35.425 0.76 ;
      LAYER metal2 ;
        RECT 36.5825 0.77 36.6525 0.905 ;
        RECT 36.41 0.77 36.6525 0.84 ;
        RECT 36.41 0.55 36.48 0.84 ;
        RECT 35.65 0.55 36.48 0.62 ;
        RECT 35.8025 0.55 35.8725 0.7 ;
        RECT 35.285 0.69 35.72 0.76 ;
        RECT 35.65 0.55 35.72 0.76 ;
      LAYER metal1 ;
        RECT 36.585 0.77 36.65 0.905 ;
        RECT 35.805 0.565 35.87 0.7 ;
        RECT 35.285 0.6925 35.42 0.7575 ;
        RECT 35.285 0.69 35.35 0.825 ;
      LAYER via2 ;
        RECT 35.32 0.69 35.39 0.76 ;
      LAYER via1 ;
        RECT 35.32 0.6925 35.385 0.7575 ;
        RECT 35.805 0.6 35.87 0.665 ;
        RECT 36.585 0.805 36.65 0.87 ;
    END
  END rd_sel[18]
  PIN rd_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 32.585 0.69 32.725 0.76 ;
      LAYER metal2 ;
        RECT 33.8825 0.77 33.9525 0.905 ;
        RECT 33.71 0.77 33.9525 0.84 ;
        RECT 33.71 0.55 33.78 0.84 ;
        RECT 32.95 0.55 33.78 0.62 ;
        RECT 33.1025 0.55 33.1725 0.7 ;
        RECT 32.585 0.69 33.02 0.76 ;
        RECT 32.95 0.55 33.02 0.76 ;
      LAYER metal1 ;
        RECT 33.885 0.77 33.95 0.905 ;
        RECT 33.105 0.565 33.17 0.7 ;
        RECT 32.585 0.6925 32.72 0.7575 ;
        RECT 32.585 0.69 32.65 0.825 ;
      LAYER via2 ;
        RECT 32.62 0.69 32.69 0.76 ;
      LAYER via1 ;
        RECT 32.62 0.6925 32.685 0.7575 ;
        RECT 33.105 0.6 33.17 0.665 ;
        RECT 33.885 0.805 33.95 0.87 ;
    END
  END rd_sel[19]
  PIN rd_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 81.185 0.69 81.325 0.76 ;
      LAYER metal2 ;
        RECT 82.4825 0.77 82.5525 0.905 ;
        RECT 82.31 0.77 82.5525 0.84 ;
        RECT 82.31 0.55 82.38 0.84 ;
        RECT 81.55 0.55 82.38 0.62 ;
        RECT 81.7025 0.55 81.7725 0.7 ;
        RECT 81.185 0.69 81.62 0.76 ;
        RECT 81.55 0.55 81.62 0.76 ;
      LAYER metal1 ;
        RECT 82.485 0.77 82.55 0.905 ;
        RECT 81.705 0.565 81.77 0.7 ;
        RECT 81.185 0.6925 81.32 0.7575 ;
        RECT 81.185 0.69 81.25 0.825 ;
      LAYER via2 ;
        RECT 81.22 0.69 81.29 0.76 ;
      LAYER via1 ;
        RECT 81.22 0.6925 81.285 0.7575 ;
        RECT 81.705 0.6 81.77 0.665 ;
        RECT 82.485 0.805 82.55 0.87 ;
    END
  END rd_sel[1]
  PIN rd_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 29.885 0.69 30.025 0.76 ;
      LAYER metal2 ;
        RECT 31.1825 0.77 31.2525 0.905 ;
        RECT 31.01 0.77 31.2525 0.84 ;
        RECT 31.01 0.55 31.08 0.84 ;
        RECT 30.25 0.55 31.08 0.62 ;
        RECT 30.4025 0.55 30.4725 0.7 ;
        RECT 29.885 0.69 30.32 0.76 ;
        RECT 30.25 0.55 30.32 0.76 ;
      LAYER metal1 ;
        RECT 31.185 0.77 31.25 0.905 ;
        RECT 30.405 0.565 30.47 0.7 ;
        RECT 29.885 0.6925 30.02 0.7575 ;
        RECT 29.885 0.69 29.95 0.825 ;
      LAYER via2 ;
        RECT 29.92 0.69 29.99 0.76 ;
      LAYER via1 ;
        RECT 29.92 0.6925 29.985 0.7575 ;
        RECT 30.405 0.6 30.47 0.665 ;
        RECT 31.185 0.805 31.25 0.87 ;
    END
  END rd_sel[20]
  PIN rd_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 27.185 0.69 27.325 0.76 ;
      LAYER metal2 ;
        RECT 28.4825 0.77 28.5525 0.905 ;
        RECT 28.31 0.77 28.5525 0.84 ;
        RECT 28.31 0.55 28.38 0.84 ;
        RECT 27.55 0.55 28.38 0.62 ;
        RECT 27.7025 0.55 27.7725 0.7 ;
        RECT 27.185 0.69 27.62 0.76 ;
        RECT 27.55 0.55 27.62 0.76 ;
      LAYER metal1 ;
        RECT 28.485 0.77 28.55 0.905 ;
        RECT 27.705 0.565 27.77 0.7 ;
        RECT 27.185 0.6925 27.32 0.7575 ;
        RECT 27.185 0.69 27.25 0.825 ;
      LAYER via2 ;
        RECT 27.22 0.69 27.29 0.76 ;
      LAYER via1 ;
        RECT 27.22 0.6925 27.285 0.7575 ;
        RECT 27.705 0.6 27.77 0.665 ;
        RECT 28.485 0.805 28.55 0.87 ;
    END
  END rd_sel[21]
  PIN rd_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 24.485 0.69 24.625 0.76 ;
      LAYER metal2 ;
        RECT 25.7825 0.77 25.8525 0.905 ;
        RECT 25.61 0.77 25.8525 0.84 ;
        RECT 25.61 0.55 25.68 0.84 ;
        RECT 24.85 0.55 25.68 0.62 ;
        RECT 25.0025 0.55 25.0725 0.7 ;
        RECT 24.485 0.69 24.92 0.76 ;
        RECT 24.85 0.55 24.92 0.76 ;
      LAYER metal1 ;
        RECT 25.785 0.77 25.85 0.905 ;
        RECT 25.005 0.565 25.07 0.7 ;
        RECT 24.485 0.6925 24.62 0.7575 ;
        RECT 24.485 0.69 24.55 0.825 ;
      LAYER via2 ;
        RECT 24.52 0.69 24.59 0.76 ;
      LAYER via1 ;
        RECT 24.52 0.6925 24.585 0.7575 ;
        RECT 25.005 0.6 25.07 0.665 ;
        RECT 25.785 0.805 25.85 0.87 ;
    END
  END rd_sel[22]
  PIN rd_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 21.785 0.69 21.925 0.76 ;
      LAYER metal2 ;
        RECT 23.0825 0.77 23.1525 0.905 ;
        RECT 22.91 0.77 23.1525 0.84 ;
        RECT 22.91 0.55 22.98 0.84 ;
        RECT 22.15 0.55 22.98 0.62 ;
        RECT 22.3025 0.55 22.3725 0.7 ;
        RECT 21.785 0.69 22.22 0.76 ;
        RECT 22.15 0.55 22.22 0.76 ;
      LAYER metal1 ;
        RECT 23.085 0.77 23.15 0.905 ;
        RECT 22.305 0.565 22.37 0.7 ;
        RECT 21.785 0.6925 21.92 0.7575 ;
        RECT 21.785 0.69 21.85 0.825 ;
      LAYER via2 ;
        RECT 21.82 0.69 21.89 0.76 ;
      LAYER via1 ;
        RECT 21.82 0.6925 21.885 0.7575 ;
        RECT 22.305 0.6 22.37 0.665 ;
        RECT 23.085 0.805 23.15 0.87 ;
    END
  END rd_sel[23]
  PIN rd_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 19.085 0.69 19.225 0.76 ;
      LAYER metal2 ;
        RECT 20.3825 0.77 20.4525 0.905 ;
        RECT 20.21 0.77 20.4525 0.84 ;
        RECT 20.21 0.55 20.28 0.84 ;
        RECT 19.45 0.55 20.28 0.62 ;
        RECT 19.6025 0.55 19.6725 0.7 ;
        RECT 19.085 0.69 19.52 0.76 ;
        RECT 19.45 0.55 19.52 0.76 ;
      LAYER metal1 ;
        RECT 20.385 0.77 20.45 0.905 ;
        RECT 19.605 0.565 19.67 0.7 ;
        RECT 19.085 0.6925 19.22 0.7575 ;
        RECT 19.085 0.69 19.15 0.825 ;
      LAYER via2 ;
        RECT 19.12 0.69 19.19 0.76 ;
      LAYER via1 ;
        RECT 19.12 0.6925 19.185 0.7575 ;
        RECT 19.605 0.6 19.67 0.665 ;
        RECT 20.385 0.805 20.45 0.87 ;
    END
  END rd_sel[24]
  PIN rd_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 16.385 0.69 16.525 0.76 ;
      LAYER metal2 ;
        RECT 17.6825 0.77 17.7525 0.905 ;
        RECT 17.51 0.77 17.7525 0.84 ;
        RECT 17.51 0.55 17.58 0.84 ;
        RECT 16.75 0.55 17.58 0.62 ;
        RECT 16.9025 0.55 16.9725 0.7 ;
        RECT 16.385 0.69 16.82 0.76 ;
        RECT 16.75 0.55 16.82 0.76 ;
      LAYER metal1 ;
        RECT 17.685 0.77 17.75 0.905 ;
        RECT 16.905 0.565 16.97 0.7 ;
        RECT 16.385 0.6925 16.52 0.7575 ;
        RECT 16.385 0.69 16.45 0.825 ;
      LAYER via2 ;
        RECT 16.42 0.69 16.49 0.76 ;
      LAYER via1 ;
        RECT 16.42 0.6925 16.485 0.7575 ;
        RECT 16.905 0.6 16.97 0.665 ;
        RECT 17.685 0.805 17.75 0.87 ;
    END
  END rd_sel[25]
  PIN rd_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 13.685 0.69 13.825 0.76 ;
      LAYER metal2 ;
        RECT 14.9825 0.77 15.0525 0.905 ;
        RECT 14.81 0.77 15.0525 0.84 ;
        RECT 14.81 0.55 14.88 0.84 ;
        RECT 14.05 0.55 14.88 0.62 ;
        RECT 14.2025 0.55 14.2725 0.7 ;
        RECT 13.685 0.69 14.12 0.76 ;
        RECT 14.05 0.55 14.12 0.76 ;
      LAYER metal1 ;
        RECT 14.985 0.77 15.05 0.905 ;
        RECT 14.205 0.565 14.27 0.7 ;
        RECT 13.685 0.6925 13.82 0.7575 ;
        RECT 13.685 0.69 13.75 0.825 ;
      LAYER via2 ;
        RECT 13.72 0.69 13.79 0.76 ;
      LAYER via1 ;
        RECT 13.72 0.6925 13.785 0.7575 ;
        RECT 14.205 0.6 14.27 0.665 ;
        RECT 14.985 0.805 15.05 0.87 ;
    END
  END rd_sel[26]
  PIN rd_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 10.985 0.69 11.125 0.76 ;
      LAYER metal2 ;
        RECT 12.2825 0.77 12.3525 0.905 ;
        RECT 12.11 0.77 12.3525 0.84 ;
        RECT 12.11 0.55 12.18 0.84 ;
        RECT 11.35 0.55 12.18 0.62 ;
        RECT 11.5025 0.55 11.5725 0.7 ;
        RECT 10.985 0.69 11.42 0.76 ;
        RECT 11.35 0.55 11.42 0.76 ;
      LAYER metal1 ;
        RECT 12.285 0.77 12.35 0.905 ;
        RECT 11.505 0.565 11.57 0.7 ;
        RECT 10.985 0.6925 11.12 0.7575 ;
        RECT 10.985 0.69 11.05 0.825 ;
      LAYER via2 ;
        RECT 11.02 0.69 11.09 0.76 ;
      LAYER via1 ;
        RECT 11.02 0.6925 11.085 0.7575 ;
        RECT 11.505 0.6 11.57 0.665 ;
        RECT 12.285 0.805 12.35 0.87 ;
    END
  END rd_sel[27]
  PIN rd_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 8.285 0.69 8.425 0.76 ;
      LAYER metal2 ;
        RECT 9.5825 0.77 9.6525 0.905 ;
        RECT 9.41 0.77 9.6525 0.84 ;
        RECT 9.41 0.55 9.48 0.84 ;
        RECT 8.65 0.55 9.48 0.62 ;
        RECT 8.8025 0.55 8.8725 0.7 ;
        RECT 8.285 0.69 8.72 0.76 ;
        RECT 8.65 0.55 8.72 0.76 ;
      LAYER metal1 ;
        RECT 9.585 0.77 9.65 0.905 ;
        RECT 8.805 0.565 8.87 0.7 ;
        RECT 8.285 0.6925 8.42 0.7575 ;
        RECT 8.285 0.69 8.35 0.825 ;
      LAYER via2 ;
        RECT 8.32 0.69 8.39 0.76 ;
      LAYER via1 ;
        RECT 8.32 0.6925 8.385 0.7575 ;
        RECT 8.805 0.6 8.87 0.665 ;
        RECT 9.585 0.805 9.65 0.87 ;
    END
  END rd_sel[28]
  PIN rd_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 5.585 0.69 5.725 0.76 ;
      LAYER metal2 ;
        RECT 6.8825 0.77 6.9525 0.905 ;
        RECT 6.71 0.77 6.9525 0.84 ;
        RECT 6.71 0.55 6.78 0.84 ;
        RECT 5.95 0.55 6.78 0.62 ;
        RECT 6.1025 0.55 6.1725 0.7 ;
        RECT 5.585 0.69 6.02 0.76 ;
        RECT 5.95 0.55 6.02 0.76 ;
      LAYER metal1 ;
        RECT 6.885 0.77 6.95 0.905 ;
        RECT 6.105 0.565 6.17 0.7 ;
        RECT 5.585 0.6925 5.72 0.7575 ;
        RECT 5.585 0.69 5.65 0.825 ;
      LAYER via2 ;
        RECT 5.62 0.69 5.69 0.76 ;
      LAYER via1 ;
        RECT 5.62 0.6925 5.685 0.7575 ;
        RECT 6.105 0.6 6.17 0.665 ;
        RECT 6.885 0.805 6.95 0.87 ;
    END
  END rd_sel[29]
  PIN rd_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 78.485 0.69 78.625 0.76 ;
      LAYER metal2 ;
        RECT 79.7825 0.77 79.8525 0.905 ;
        RECT 79.61 0.77 79.8525 0.84 ;
        RECT 79.61 0.55 79.68 0.84 ;
        RECT 78.85 0.55 79.68 0.62 ;
        RECT 79.0025 0.55 79.0725 0.7 ;
        RECT 78.485 0.69 78.92 0.76 ;
        RECT 78.85 0.55 78.92 0.76 ;
      LAYER metal1 ;
        RECT 79.785 0.77 79.85 0.905 ;
        RECT 79.005 0.565 79.07 0.7 ;
        RECT 78.485 0.6925 78.62 0.7575 ;
        RECT 78.485 0.69 78.55 0.825 ;
      LAYER via2 ;
        RECT 78.52 0.69 78.59 0.76 ;
      LAYER via1 ;
        RECT 78.52 0.6925 78.585 0.7575 ;
        RECT 79.005 0.6 79.07 0.665 ;
        RECT 79.785 0.805 79.85 0.87 ;
    END
  END rd_sel[2]
  PIN rd_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 2.885 0.69 3.025 0.76 ;
      LAYER metal2 ;
        RECT 4.1825 0.77 4.2525 0.905 ;
        RECT 4.01 0.77 4.2525 0.84 ;
        RECT 4.01 0.55 4.08 0.84 ;
        RECT 3.25 0.55 4.08 0.62 ;
        RECT 3.4025 0.55 3.4725 0.7 ;
        RECT 2.885 0.69 3.32 0.76 ;
        RECT 3.25 0.55 3.32 0.76 ;
      LAYER metal1 ;
        RECT 4.185 0.77 4.25 0.905 ;
        RECT 3.405 0.565 3.47 0.7 ;
        RECT 2.885 0.6925 3.02 0.7575 ;
        RECT 2.885 0.69 2.95 0.825 ;
      LAYER via2 ;
        RECT 2.92 0.69 2.99 0.76 ;
      LAYER via1 ;
        RECT 2.92 0.6925 2.985 0.7575 ;
        RECT 3.405 0.6 3.47 0.665 ;
        RECT 4.185 0.805 4.25 0.87 ;
    END
  END rd_sel[30]
  PIN rd_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.185 0.69 0.325 0.76 ;
      LAYER metal2 ;
        RECT 1.4825 0.77 1.5525 0.905 ;
        RECT 1.31 0.77 1.5525 0.84 ;
        RECT 1.31 0.55 1.38 0.84 ;
        RECT 0.55 0.55 1.38 0.62 ;
        RECT 0.7025 0.55 0.7725 0.7 ;
        RECT 0.185 0.69 0.62 0.76 ;
        RECT 0.55 0.55 0.62 0.76 ;
      LAYER metal1 ;
        RECT 1.485 0.77 1.55 0.905 ;
        RECT 0.705 0.565 0.77 0.7 ;
        RECT 0.185 0.6925 0.32 0.7575 ;
        RECT 0.185 0.69 0.25 0.825 ;
      LAYER via2 ;
        RECT 0.22 0.69 0.29 0.76 ;
      LAYER via1 ;
        RECT 0.22 0.6925 0.285 0.7575 ;
        RECT 0.705 0.6 0.77 0.665 ;
        RECT 1.485 0.805 1.55 0.87 ;
    END
  END rd_sel[31]
  PIN rd_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.785 0.69 75.925 0.76 ;
      LAYER metal2 ;
        RECT 77.0825 0.77 77.1525 0.905 ;
        RECT 76.91 0.77 77.1525 0.84 ;
        RECT 76.91 0.55 76.98 0.84 ;
        RECT 76.15 0.55 76.98 0.62 ;
        RECT 76.3025 0.55 76.3725 0.7 ;
        RECT 75.785 0.69 76.22 0.76 ;
        RECT 76.15 0.55 76.22 0.76 ;
      LAYER metal1 ;
        RECT 77.085 0.77 77.15 0.905 ;
        RECT 76.305 0.565 76.37 0.7 ;
        RECT 75.785 0.6925 75.92 0.7575 ;
        RECT 75.785 0.69 75.85 0.825 ;
      LAYER via2 ;
        RECT 75.82 0.69 75.89 0.76 ;
      LAYER via1 ;
        RECT 75.82 0.6925 75.885 0.7575 ;
        RECT 76.305 0.6 76.37 0.665 ;
        RECT 77.085 0.805 77.15 0.87 ;
    END
  END rd_sel[3]
  PIN rd_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 73.085 0.69 73.225 0.76 ;
      LAYER metal2 ;
        RECT 74.3825 0.77 74.4525 0.905 ;
        RECT 74.21 0.77 74.4525 0.84 ;
        RECT 74.21 0.55 74.28 0.84 ;
        RECT 73.45 0.55 74.28 0.62 ;
        RECT 73.6025 0.55 73.6725 0.7 ;
        RECT 73.085 0.69 73.52 0.76 ;
        RECT 73.45 0.55 73.52 0.76 ;
      LAYER metal1 ;
        RECT 74.385 0.77 74.45 0.905 ;
        RECT 73.605 0.565 73.67 0.7 ;
        RECT 73.085 0.6925 73.22 0.7575 ;
        RECT 73.085 0.69 73.15 0.825 ;
      LAYER via2 ;
        RECT 73.12 0.69 73.19 0.76 ;
      LAYER via1 ;
        RECT 73.12 0.6925 73.185 0.7575 ;
        RECT 73.605 0.6 73.67 0.665 ;
        RECT 74.385 0.805 74.45 0.87 ;
    END
  END rd_sel[4]
  PIN rd_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 70.385 0.69 70.525 0.76 ;
      LAYER metal2 ;
        RECT 71.6825 0.77 71.7525 0.905 ;
        RECT 71.51 0.77 71.7525 0.84 ;
        RECT 71.51 0.55 71.58 0.84 ;
        RECT 70.75 0.55 71.58 0.62 ;
        RECT 70.9025 0.55 70.9725 0.7 ;
        RECT 70.385 0.69 70.82 0.76 ;
        RECT 70.75 0.55 70.82 0.76 ;
      LAYER metal1 ;
        RECT 71.685 0.77 71.75 0.905 ;
        RECT 70.905 0.565 70.97 0.7 ;
        RECT 70.385 0.6925 70.52 0.7575 ;
        RECT 70.385 0.69 70.45 0.825 ;
      LAYER via2 ;
        RECT 70.42 0.69 70.49 0.76 ;
      LAYER via1 ;
        RECT 70.42 0.6925 70.485 0.7575 ;
        RECT 70.905 0.6 70.97 0.665 ;
        RECT 71.685 0.805 71.75 0.87 ;
    END
  END rd_sel[5]
  PIN rd_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 67.685 0.69 67.825 0.76 ;
      LAYER metal2 ;
        RECT 68.9825 0.77 69.0525 0.905 ;
        RECT 68.81 0.77 69.0525 0.84 ;
        RECT 68.81 0.55 68.88 0.84 ;
        RECT 68.05 0.55 68.88 0.62 ;
        RECT 68.2025 0.55 68.2725 0.7 ;
        RECT 67.685 0.69 68.12 0.76 ;
        RECT 68.05 0.55 68.12 0.76 ;
      LAYER metal1 ;
        RECT 68.985 0.77 69.05 0.905 ;
        RECT 68.205 0.565 68.27 0.7 ;
        RECT 67.685 0.6925 67.82 0.7575 ;
        RECT 67.685 0.69 67.75 0.825 ;
      LAYER via2 ;
        RECT 67.72 0.69 67.79 0.76 ;
      LAYER via1 ;
        RECT 67.72 0.6925 67.785 0.7575 ;
        RECT 68.205 0.6 68.27 0.665 ;
        RECT 68.985 0.805 69.05 0.87 ;
    END
  END rd_sel[6]
  PIN rd_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 64.985 0.69 65.125 0.76 ;
      LAYER metal2 ;
        RECT 66.2825 0.77 66.3525 0.905 ;
        RECT 66.11 0.77 66.3525 0.84 ;
        RECT 66.11 0.55 66.18 0.84 ;
        RECT 65.35 0.55 66.18 0.62 ;
        RECT 65.5025 0.55 65.5725 0.7 ;
        RECT 64.985 0.69 65.42 0.76 ;
        RECT 65.35 0.55 65.42 0.76 ;
      LAYER metal1 ;
        RECT 66.285 0.77 66.35 0.905 ;
        RECT 65.505 0.565 65.57 0.7 ;
        RECT 64.985 0.6925 65.12 0.7575 ;
        RECT 64.985 0.69 65.05 0.825 ;
      LAYER via2 ;
        RECT 65.02 0.69 65.09 0.76 ;
      LAYER via1 ;
        RECT 65.02 0.6925 65.085 0.7575 ;
        RECT 65.505 0.6 65.57 0.665 ;
        RECT 66.285 0.805 66.35 0.87 ;
    END
  END rd_sel[7]
  PIN rd_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 62.285 0.69 62.425 0.76 ;
      LAYER metal2 ;
        RECT 63.5825 0.77 63.6525 0.905 ;
        RECT 63.41 0.77 63.6525 0.84 ;
        RECT 63.41 0.55 63.48 0.84 ;
        RECT 62.65 0.55 63.48 0.62 ;
        RECT 62.8025 0.55 62.8725 0.7 ;
        RECT 62.285 0.69 62.72 0.76 ;
        RECT 62.65 0.55 62.72 0.76 ;
      LAYER metal1 ;
        RECT 63.585 0.77 63.65 0.905 ;
        RECT 62.805 0.565 62.87 0.7 ;
        RECT 62.285 0.6925 62.42 0.7575 ;
        RECT 62.285 0.69 62.35 0.825 ;
      LAYER via2 ;
        RECT 62.32 0.69 62.39 0.76 ;
      LAYER via1 ;
        RECT 62.32 0.6925 62.385 0.7575 ;
        RECT 62.805 0.6 62.87 0.665 ;
        RECT 63.585 0.805 63.65 0.87 ;
    END
  END rd_sel[8]
  PIN rd_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 59.585 0.69 59.725 0.76 ;
      LAYER metal2 ;
        RECT 60.8825 0.77 60.9525 0.905 ;
        RECT 60.71 0.77 60.9525 0.84 ;
        RECT 60.71 0.55 60.78 0.84 ;
        RECT 59.95 0.55 60.78 0.62 ;
        RECT 60.1025 0.55 60.1725 0.7 ;
        RECT 59.585 0.69 60.02 0.76 ;
        RECT 59.95 0.55 60.02 0.76 ;
      LAYER metal1 ;
        RECT 60.885 0.77 60.95 0.905 ;
        RECT 60.105 0.565 60.17 0.7 ;
        RECT 59.585 0.6925 59.72 0.7575 ;
        RECT 59.585 0.69 59.65 0.825 ;
      LAYER via2 ;
        RECT 59.62 0.69 59.69 0.76 ;
      LAYER via1 ;
        RECT 59.62 0.6925 59.685 0.7575 ;
        RECT 60.105 0.6 60.17 0.665 ;
        RECT 60.885 0.805 60.95 0.87 ;
    END
  END rd_sel[9]
  PIN rs1_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 86.28 0.69 86.345 0.825 ;
        RECT 86.05 0.725 86.345 0.79 ;
        RECT 86.05 0.265 86.115 1.14 ;
    END
  END rs1_rdata
  PIN rs1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.4025 0.41 84.4725 0.545 ;
        RECT 83.995 0.41 84.4725 0.48 ;
        RECT 83.93 0.52 84.065 0.59 ;
        RECT 83.995 0.41 84.065 0.59 ;
      LAYER metal1 ;
        RECT 84.405 0.41 84.47 0.545 ;
        RECT 83.93 0.5225 84.065 0.5875 ;
        RECT 83.995 0.49 84.06 0.625 ;
      LAYER via1 ;
        RECT 83.965 0.5225 84.03 0.5875 ;
        RECT 84.405 0.445 84.47 0.51 ;
    END
  END rs1_sel[0]
  PIN rs1_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 56.9225 0.535 57.0625 0.605 ;
      LAYER metal2 ;
        RECT 58.5875 0.41 58.6575 0.545 ;
        RECT 56.9925 0.41 58.6575 0.48 ;
        RECT 56.9225 0.535 57.0625 0.605 ;
        RECT 56.9925 0.41 57.0625 0.605 ;
      LAYER metal1 ;
        RECT 58.59 0.41 58.655 0.545 ;
        RECT 56.9275 0.5375 57.0625 0.6025 ;
        RECT 56.995 0.49 57.06 0.625 ;
      LAYER via2 ;
        RECT 56.9575 0.535 57.0275 0.605 ;
      LAYER via1 ;
        RECT 56.9625 0.5375 57.0275 0.6025 ;
        RECT 58.59 0.445 58.655 0.51 ;
    END
  END rs1_sel[10]
  PIN rs1_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 54.2225 0.535 54.3625 0.605 ;
      LAYER metal2 ;
        RECT 55.8875 0.41 55.9575 0.545 ;
        RECT 54.2925 0.41 55.9575 0.48 ;
        RECT 54.2225 0.535 54.3625 0.605 ;
        RECT 54.2925 0.41 54.3625 0.605 ;
      LAYER metal1 ;
        RECT 55.89 0.41 55.955 0.545 ;
        RECT 54.2275 0.5375 54.3625 0.6025 ;
        RECT 54.295 0.49 54.36 0.625 ;
      LAYER via2 ;
        RECT 54.2575 0.535 54.3275 0.605 ;
      LAYER via1 ;
        RECT 54.2625 0.5375 54.3275 0.6025 ;
        RECT 55.89 0.445 55.955 0.51 ;
    END
  END rs1_sel[11]
  PIN rs1_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 51.5225 0.535 51.6625 0.605 ;
      LAYER metal2 ;
        RECT 53.1875 0.41 53.2575 0.545 ;
        RECT 51.5925 0.41 53.2575 0.48 ;
        RECT 51.5225 0.535 51.6625 0.605 ;
        RECT 51.5925 0.41 51.6625 0.605 ;
      LAYER metal1 ;
        RECT 53.19 0.41 53.255 0.545 ;
        RECT 51.5275 0.5375 51.6625 0.6025 ;
        RECT 51.595 0.49 51.66 0.625 ;
      LAYER via2 ;
        RECT 51.5575 0.535 51.6275 0.605 ;
      LAYER via1 ;
        RECT 51.5625 0.5375 51.6275 0.6025 ;
        RECT 53.19 0.445 53.255 0.51 ;
    END
  END rs1_sel[12]
  PIN rs1_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 48.8225 0.535 48.9625 0.605 ;
      LAYER metal2 ;
        RECT 50.4875 0.41 50.5575 0.545 ;
        RECT 48.8925 0.41 50.5575 0.48 ;
        RECT 48.8225 0.535 48.9625 0.605 ;
        RECT 48.8925 0.41 48.9625 0.605 ;
      LAYER metal1 ;
        RECT 50.49 0.41 50.555 0.545 ;
        RECT 48.8275 0.5375 48.9625 0.6025 ;
        RECT 48.895 0.49 48.96 0.625 ;
      LAYER via2 ;
        RECT 48.8575 0.535 48.9275 0.605 ;
      LAYER via1 ;
        RECT 48.8625 0.5375 48.9275 0.6025 ;
        RECT 50.49 0.445 50.555 0.51 ;
    END
  END rs1_sel[13]
  PIN rs1_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 46.1225 0.535 46.2625 0.605 ;
      LAYER metal2 ;
        RECT 47.7875 0.41 47.8575 0.545 ;
        RECT 46.1925 0.41 47.8575 0.48 ;
        RECT 46.1225 0.535 46.2625 0.605 ;
        RECT 46.1925 0.41 46.2625 0.605 ;
      LAYER metal1 ;
        RECT 47.79 0.41 47.855 0.545 ;
        RECT 46.1275 0.5375 46.2625 0.6025 ;
        RECT 46.195 0.49 46.26 0.625 ;
      LAYER via2 ;
        RECT 46.1575 0.535 46.2275 0.605 ;
      LAYER via1 ;
        RECT 46.1625 0.5375 46.2275 0.6025 ;
        RECT 47.79 0.445 47.855 0.51 ;
    END
  END rs1_sel[14]
  PIN rs1_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 43.4225 0.535 43.5625 0.605 ;
      LAYER metal2 ;
        RECT 45.0875 0.41 45.1575 0.545 ;
        RECT 43.4925 0.41 45.1575 0.48 ;
        RECT 43.4225 0.535 43.5625 0.605 ;
        RECT 43.4925 0.41 43.5625 0.605 ;
      LAYER metal1 ;
        RECT 45.09 0.41 45.155 0.545 ;
        RECT 43.4275 0.5375 43.5625 0.6025 ;
        RECT 43.495 0.49 43.56 0.625 ;
      LAYER via2 ;
        RECT 43.4575 0.535 43.5275 0.605 ;
      LAYER via1 ;
        RECT 43.4625 0.5375 43.5275 0.6025 ;
        RECT 45.09 0.445 45.155 0.51 ;
    END
  END rs1_sel[15]
  PIN rs1_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 40.7225 0.535 40.8625 0.605 ;
      LAYER metal2 ;
        RECT 42.3875 0.41 42.4575 0.545 ;
        RECT 40.7925 0.41 42.4575 0.48 ;
        RECT 40.7225 0.535 40.8625 0.605 ;
        RECT 40.7925 0.41 40.8625 0.605 ;
      LAYER metal1 ;
        RECT 42.39 0.41 42.455 0.545 ;
        RECT 40.7275 0.5375 40.8625 0.6025 ;
        RECT 40.795 0.49 40.86 0.625 ;
      LAYER via2 ;
        RECT 40.7575 0.535 40.8275 0.605 ;
      LAYER via1 ;
        RECT 40.7625 0.5375 40.8275 0.6025 ;
        RECT 42.39 0.445 42.455 0.51 ;
    END
  END rs1_sel[16]
  PIN rs1_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 38.0225 0.535 38.1625 0.605 ;
      LAYER metal2 ;
        RECT 39.6875 0.41 39.7575 0.545 ;
        RECT 38.0925 0.41 39.7575 0.48 ;
        RECT 38.0225 0.535 38.1625 0.605 ;
        RECT 38.0925 0.41 38.1625 0.605 ;
      LAYER metal1 ;
        RECT 39.69 0.41 39.755 0.545 ;
        RECT 38.0275 0.5375 38.1625 0.6025 ;
        RECT 38.095 0.49 38.16 0.625 ;
      LAYER via2 ;
        RECT 38.0575 0.535 38.1275 0.605 ;
      LAYER via1 ;
        RECT 38.0625 0.5375 38.1275 0.6025 ;
        RECT 39.69 0.445 39.755 0.51 ;
    END
  END rs1_sel[17]
  PIN rs1_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 35.3225 0.535 35.4625 0.605 ;
      LAYER metal2 ;
        RECT 36.9875 0.41 37.0575 0.545 ;
        RECT 35.3925 0.41 37.0575 0.48 ;
        RECT 35.3225 0.535 35.4625 0.605 ;
        RECT 35.3925 0.41 35.4625 0.605 ;
      LAYER metal1 ;
        RECT 36.99 0.41 37.055 0.545 ;
        RECT 35.3275 0.5375 35.4625 0.6025 ;
        RECT 35.395 0.49 35.46 0.625 ;
      LAYER via2 ;
        RECT 35.3575 0.535 35.4275 0.605 ;
      LAYER via1 ;
        RECT 35.3625 0.5375 35.4275 0.6025 ;
        RECT 36.99 0.445 37.055 0.51 ;
    END
  END rs1_sel[18]
  PIN rs1_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 32.6225 0.535 32.7625 0.605 ;
      LAYER metal2 ;
        RECT 34.2875 0.41 34.3575 0.545 ;
        RECT 32.6925 0.41 34.3575 0.48 ;
        RECT 32.6225 0.535 32.7625 0.605 ;
        RECT 32.6925 0.41 32.7625 0.605 ;
      LAYER metal1 ;
        RECT 34.29 0.41 34.355 0.545 ;
        RECT 32.6275 0.5375 32.7625 0.6025 ;
        RECT 32.695 0.49 32.76 0.625 ;
      LAYER via2 ;
        RECT 32.6575 0.535 32.7275 0.605 ;
      LAYER via1 ;
        RECT 32.6625 0.5375 32.7275 0.6025 ;
        RECT 34.29 0.445 34.355 0.51 ;
    END
  END rs1_sel[19]
  PIN rs1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 81.2225 0.535 81.3625 0.605 ;
      LAYER metal2 ;
        RECT 82.8875 0.41 82.9575 0.545 ;
        RECT 81.2925 0.41 82.9575 0.48 ;
        RECT 81.2225 0.535 81.3625 0.605 ;
        RECT 81.2925 0.41 81.3625 0.605 ;
      LAYER metal1 ;
        RECT 82.89 0.41 82.955 0.545 ;
        RECT 81.2275 0.5375 81.3625 0.6025 ;
        RECT 81.295 0.49 81.36 0.625 ;
      LAYER via2 ;
        RECT 81.2575 0.535 81.3275 0.605 ;
      LAYER via1 ;
        RECT 81.2625 0.5375 81.3275 0.6025 ;
        RECT 82.89 0.445 82.955 0.51 ;
    END
  END rs1_sel[1]
  PIN rs1_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 29.9225 0.535 30.0625 0.605 ;
      LAYER metal2 ;
        RECT 31.5875 0.41 31.6575 0.545 ;
        RECT 29.9925 0.41 31.6575 0.48 ;
        RECT 29.9225 0.535 30.0625 0.605 ;
        RECT 29.9925 0.41 30.0625 0.605 ;
      LAYER metal1 ;
        RECT 31.59 0.41 31.655 0.545 ;
        RECT 29.9275 0.5375 30.0625 0.6025 ;
        RECT 29.995 0.49 30.06 0.625 ;
      LAYER via2 ;
        RECT 29.9575 0.535 30.0275 0.605 ;
      LAYER via1 ;
        RECT 29.9625 0.5375 30.0275 0.6025 ;
        RECT 31.59 0.445 31.655 0.51 ;
    END
  END rs1_sel[20]
  PIN rs1_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 27.2225 0.535 27.3625 0.605 ;
      LAYER metal2 ;
        RECT 28.8875 0.41 28.9575 0.545 ;
        RECT 27.2925 0.41 28.9575 0.48 ;
        RECT 27.2225 0.535 27.3625 0.605 ;
        RECT 27.2925 0.41 27.3625 0.605 ;
      LAYER metal1 ;
        RECT 28.89 0.41 28.955 0.545 ;
        RECT 27.2275 0.5375 27.3625 0.6025 ;
        RECT 27.295 0.49 27.36 0.625 ;
      LAYER via2 ;
        RECT 27.2575 0.535 27.3275 0.605 ;
      LAYER via1 ;
        RECT 27.2625 0.5375 27.3275 0.6025 ;
        RECT 28.89 0.445 28.955 0.51 ;
    END
  END rs1_sel[21]
  PIN rs1_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 24.5225 0.535 24.6625 0.605 ;
      LAYER metal2 ;
        RECT 26.1875 0.41 26.2575 0.545 ;
        RECT 24.5925 0.41 26.2575 0.48 ;
        RECT 24.5225 0.535 24.6625 0.605 ;
        RECT 24.5925 0.41 24.6625 0.605 ;
      LAYER metal1 ;
        RECT 26.19 0.41 26.255 0.545 ;
        RECT 24.5275 0.5375 24.6625 0.6025 ;
        RECT 24.595 0.49 24.66 0.625 ;
      LAYER via2 ;
        RECT 24.5575 0.535 24.6275 0.605 ;
      LAYER via1 ;
        RECT 24.5625 0.5375 24.6275 0.6025 ;
        RECT 26.19 0.445 26.255 0.51 ;
    END
  END rs1_sel[22]
  PIN rs1_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 21.8225 0.535 21.9625 0.605 ;
      LAYER metal2 ;
        RECT 23.4875 0.41 23.5575 0.545 ;
        RECT 21.8925 0.41 23.5575 0.48 ;
        RECT 21.8225 0.535 21.9625 0.605 ;
        RECT 21.8925 0.41 21.9625 0.605 ;
      LAYER metal1 ;
        RECT 23.49 0.41 23.555 0.545 ;
        RECT 21.8275 0.5375 21.9625 0.6025 ;
        RECT 21.895 0.49 21.96 0.625 ;
      LAYER via2 ;
        RECT 21.8575 0.535 21.9275 0.605 ;
      LAYER via1 ;
        RECT 21.8625 0.5375 21.9275 0.6025 ;
        RECT 23.49 0.445 23.555 0.51 ;
    END
  END rs1_sel[23]
  PIN rs1_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 19.1225 0.535 19.2625 0.605 ;
      LAYER metal2 ;
        RECT 20.7875 0.41 20.8575 0.545 ;
        RECT 19.1925 0.41 20.8575 0.48 ;
        RECT 19.1225 0.535 19.2625 0.605 ;
        RECT 19.1925 0.41 19.2625 0.605 ;
      LAYER metal1 ;
        RECT 20.79 0.41 20.855 0.545 ;
        RECT 19.1275 0.5375 19.2625 0.6025 ;
        RECT 19.195 0.49 19.26 0.625 ;
      LAYER via2 ;
        RECT 19.1575 0.535 19.2275 0.605 ;
      LAYER via1 ;
        RECT 19.1625 0.5375 19.2275 0.6025 ;
        RECT 20.79 0.445 20.855 0.51 ;
    END
  END rs1_sel[24]
  PIN rs1_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 16.4225 0.535 16.5625 0.605 ;
      LAYER metal2 ;
        RECT 18.0875 0.41 18.1575 0.545 ;
        RECT 16.4925 0.41 18.1575 0.48 ;
        RECT 16.4225 0.535 16.5625 0.605 ;
        RECT 16.4925 0.41 16.5625 0.605 ;
      LAYER metal1 ;
        RECT 18.09 0.41 18.155 0.545 ;
        RECT 16.4275 0.5375 16.5625 0.6025 ;
        RECT 16.495 0.49 16.56 0.625 ;
      LAYER via2 ;
        RECT 16.4575 0.535 16.5275 0.605 ;
      LAYER via1 ;
        RECT 16.4625 0.5375 16.5275 0.6025 ;
        RECT 18.09 0.445 18.155 0.51 ;
    END
  END rs1_sel[25]
  PIN rs1_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 13.7225 0.535 13.8625 0.605 ;
      LAYER metal2 ;
        RECT 15.3875 0.41 15.4575 0.545 ;
        RECT 13.7925 0.41 15.4575 0.48 ;
        RECT 13.7225 0.535 13.8625 0.605 ;
        RECT 13.7925 0.41 13.8625 0.605 ;
      LAYER metal1 ;
        RECT 15.39 0.41 15.455 0.545 ;
        RECT 13.7275 0.5375 13.8625 0.6025 ;
        RECT 13.795 0.49 13.86 0.625 ;
      LAYER via2 ;
        RECT 13.7575 0.535 13.8275 0.605 ;
      LAYER via1 ;
        RECT 13.7625 0.5375 13.8275 0.6025 ;
        RECT 15.39 0.445 15.455 0.51 ;
    END
  END rs1_sel[26]
  PIN rs1_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 11.0225 0.535 11.1625 0.605 ;
      LAYER metal2 ;
        RECT 12.6875 0.41 12.7575 0.545 ;
        RECT 11.0925 0.41 12.7575 0.48 ;
        RECT 11.0225 0.535 11.1625 0.605 ;
        RECT 11.0925 0.41 11.1625 0.605 ;
      LAYER metal1 ;
        RECT 12.69 0.41 12.755 0.545 ;
        RECT 11.0275 0.5375 11.1625 0.6025 ;
        RECT 11.095 0.49 11.16 0.625 ;
      LAYER via2 ;
        RECT 11.0575 0.535 11.1275 0.605 ;
      LAYER via1 ;
        RECT 11.0625 0.5375 11.1275 0.6025 ;
        RECT 12.69 0.445 12.755 0.51 ;
    END
  END rs1_sel[27]
  PIN rs1_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 8.3225 0.535 8.4625 0.605 ;
      LAYER metal2 ;
        RECT 9.9875 0.41 10.0575 0.545 ;
        RECT 8.3925 0.41 10.0575 0.48 ;
        RECT 8.3225 0.535 8.4625 0.605 ;
        RECT 8.3925 0.41 8.4625 0.605 ;
      LAYER metal1 ;
        RECT 9.99 0.41 10.055 0.545 ;
        RECT 8.3275 0.5375 8.4625 0.6025 ;
        RECT 8.395 0.49 8.46 0.625 ;
      LAYER via2 ;
        RECT 8.3575 0.535 8.4275 0.605 ;
      LAYER via1 ;
        RECT 8.3625 0.5375 8.4275 0.6025 ;
        RECT 9.99 0.445 10.055 0.51 ;
    END
  END rs1_sel[28]
  PIN rs1_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 5.6225 0.535 5.7625 0.605 ;
      LAYER metal2 ;
        RECT 7.2875 0.41 7.3575 0.545 ;
        RECT 5.6925 0.41 7.3575 0.48 ;
        RECT 5.6225 0.535 5.7625 0.605 ;
        RECT 5.6925 0.41 5.7625 0.605 ;
      LAYER metal1 ;
        RECT 7.29 0.41 7.355 0.545 ;
        RECT 5.6275 0.5375 5.7625 0.6025 ;
        RECT 5.695 0.49 5.76 0.625 ;
      LAYER via2 ;
        RECT 5.6575 0.535 5.7275 0.605 ;
      LAYER via1 ;
        RECT 5.6625 0.5375 5.7275 0.6025 ;
        RECT 7.29 0.445 7.355 0.51 ;
    END
  END rs1_sel[29]
  PIN rs1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 78.5225 0.535 78.6625 0.605 ;
      LAYER metal2 ;
        RECT 80.1875 0.41 80.2575 0.545 ;
        RECT 78.5925 0.41 80.2575 0.48 ;
        RECT 78.5225 0.535 78.6625 0.605 ;
        RECT 78.5925 0.41 78.6625 0.605 ;
      LAYER metal1 ;
        RECT 80.19 0.41 80.255 0.545 ;
        RECT 78.5275 0.5375 78.6625 0.6025 ;
        RECT 78.595 0.49 78.66 0.625 ;
      LAYER via2 ;
        RECT 78.5575 0.535 78.6275 0.605 ;
      LAYER via1 ;
        RECT 78.5625 0.5375 78.6275 0.6025 ;
        RECT 80.19 0.445 80.255 0.51 ;
    END
  END rs1_sel[2]
  PIN rs1_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 2.9225 0.535 3.0625 0.605 ;
      LAYER metal2 ;
        RECT 4.5875 0.41 4.6575 0.545 ;
        RECT 2.9925 0.41 4.6575 0.48 ;
        RECT 2.9225 0.535 3.0625 0.605 ;
        RECT 2.9925 0.41 3.0625 0.605 ;
      LAYER metal1 ;
        RECT 4.59 0.41 4.655 0.545 ;
        RECT 2.9275 0.5375 3.0625 0.6025 ;
        RECT 2.995 0.49 3.06 0.625 ;
      LAYER via2 ;
        RECT 2.9575 0.535 3.0275 0.605 ;
      LAYER via1 ;
        RECT 2.9625 0.5375 3.0275 0.6025 ;
        RECT 4.59 0.445 4.655 0.51 ;
    END
  END rs1_sel[30]
  PIN rs1_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.2225 0.535 0.3625 0.605 ;
      LAYER metal2 ;
        RECT 1.8875 0.41 1.9575 0.545 ;
        RECT 0.2925 0.41 1.9575 0.48 ;
        RECT 0.2225 0.535 0.3625 0.605 ;
        RECT 0.2925 0.41 0.3625 0.605 ;
      LAYER metal1 ;
        RECT 1.89 0.41 1.955 0.545 ;
        RECT 0.2275 0.5375 0.3625 0.6025 ;
        RECT 0.295 0.49 0.36 0.625 ;
      LAYER via2 ;
        RECT 0.2575 0.535 0.3275 0.605 ;
      LAYER via1 ;
        RECT 0.2625 0.5375 0.3275 0.6025 ;
        RECT 1.89 0.445 1.955 0.51 ;
    END
  END rs1_sel[31]
  PIN rs1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.8225 0.535 75.9625 0.605 ;
      LAYER metal2 ;
        RECT 77.4875 0.41 77.5575 0.545 ;
        RECT 75.8925 0.41 77.5575 0.48 ;
        RECT 75.8225 0.535 75.9625 0.605 ;
        RECT 75.8925 0.41 75.9625 0.605 ;
      LAYER metal1 ;
        RECT 77.49 0.41 77.555 0.545 ;
        RECT 75.8275 0.5375 75.9625 0.6025 ;
        RECT 75.895 0.49 75.96 0.625 ;
      LAYER via2 ;
        RECT 75.8575 0.535 75.9275 0.605 ;
      LAYER via1 ;
        RECT 75.8625 0.5375 75.9275 0.6025 ;
        RECT 77.49 0.445 77.555 0.51 ;
    END
  END rs1_sel[3]
  PIN rs1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 73.1225 0.535 73.2625 0.605 ;
      LAYER metal2 ;
        RECT 74.7875 0.41 74.8575 0.545 ;
        RECT 73.1925 0.41 74.8575 0.48 ;
        RECT 73.1225 0.535 73.2625 0.605 ;
        RECT 73.1925 0.41 73.2625 0.605 ;
      LAYER metal1 ;
        RECT 74.79 0.41 74.855 0.545 ;
        RECT 73.1275 0.5375 73.2625 0.6025 ;
        RECT 73.195 0.49 73.26 0.625 ;
      LAYER via2 ;
        RECT 73.1575 0.535 73.2275 0.605 ;
      LAYER via1 ;
        RECT 73.1625 0.5375 73.2275 0.6025 ;
        RECT 74.79 0.445 74.855 0.51 ;
    END
  END rs1_sel[4]
  PIN rs1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 70.4225 0.535 70.5625 0.605 ;
      LAYER metal2 ;
        RECT 72.0875 0.41 72.1575 0.545 ;
        RECT 70.4925 0.41 72.1575 0.48 ;
        RECT 70.4225 0.535 70.5625 0.605 ;
        RECT 70.4925 0.41 70.5625 0.605 ;
      LAYER metal1 ;
        RECT 72.09 0.41 72.155 0.545 ;
        RECT 70.4275 0.5375 70.5625 0.6025 ;
        RECT 70.495 0.49 70.56 0.625 ;
      LAYER via2 ;
        RECT 70.4575 0.535 70.5275 0.605 ;
      LAYER via1 ;
        RECT 70.4625 0.5375 70.5275 0.6025 ;
        RECT 72.09 0.445 72.155 0.51 ;
    END
  END rs1_sel[5]
  PIN rs1_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 67.7225 0.535 67.8625 0.605 ;
      LAYER metal2 ;
        RECT 69.3875 0.41 69.4575 0.545 ;
        RECT 67.7925 0.41 69.4575 0.48 ;
        RECT 67.7225 0.535 67.8625 0.605 ;
        RECT 67.7925 0.41 67.8625 0.605 ;
      LAYER metal1 ;
        RECT 69.39 0.41 69.455 0.545 ;
        RECT 67.7275 0.5375 67.8625 0.6025 ;
        RECT 67.795 0.49 67.86 0.625 ;
      LAYER via2 ;
        RECT 67.7575 0.535 67.8275 0.605 ;
      LAYER via1 ;
        RECT 67.7625 0.5375 67.8275 0.6025 ;
        RECT 69.39 0.445 69.455 0.51 ;
    END
  END rs1_sel[6]
  PIN rs1_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 65.0225 0.535 65.1625 0.605 ;
      LAYER metal2 ;
        RECT 66.6875 0.41 66.7575 0.545 ;
        RECT 65.0925 0.41 66.7575 0.48 ;
        RECT 65.0225 0.535 65.1625 0.605 ;
        RECT 65.0925 0.41 65.1625 0.605 ;
      LAYER metal1 ;
        RECT 66.69 0.41 66.755 0.545 ;
        RECT 65.0275 0.5375 65.1625 0.6025 ;
        RECT 65.095 0.49 65.16 0.625 ;
      LAYER via2 ;
        RECT 65.0575 0.535 65.1275 0.605 ;
      LAYER via1 ;
        RECT 65.0625 0.5375 65.1275 0.6025 ;
        RECT 66.69 0.445 66.755 0.51 ;
    END
  END rs1_sel[7]
  PIN rs1_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 62.3225 0.535 62.4625 0.605 ;
      LAYER metal2 ;
        RECT 63.9875 0.41 64.0575 0.545 ;
        RECT 62.3925 0.41 64.0575 0.48 ;
        RECT 62.3225 0.535 62.4625 0.605 ;
        RECT 62.3925 0.41 62.4625 0.605 ;
      LAYER metal1 ;
        RECT 63.99 0.41 64.055 0.545 ;
        RECT 62.3275 0.5375 62.4625 0.6025 ;
        RECT 62.395 0.49 62.46 0.625 ;
      LAYER via2 ;
        RECT 62.3575 0.535 62.4275 0.605 ;
      LAYER via1 ;
        RECT 62.3625 0.5375 62.4275 0.6025 ;
        RECT 63.99 0.445 64.055 0.51 ;
    END
  END rs1_sel[8]
  PIN rs1_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 59.6225 0.535 59.7625 0.605 ;
      LAYER metal2 ;
        RECT 61.2875 0.41 61.3575 0.545 ;
        RECT 59.6925 0.41 61.3575 0.48 ;
        RECT 59.6225 0.535 59.7625 0.605 ;
        RECT 59.6925 0.41 59.7625 0.605 ;
      LAYER metal1 ;
        RECT 61.29 0.41 61.355 0.545 ;
        RECT 59.6275 0.5375 59.7625 0.6025 ;
        RECT 59.695 0.49 59.76 0.625 ;
      LAYER via2 ;
        RECT 59.6575 0.535 59.7275 0.605 ;
      LAYER via1 ;
        RECT 59.6625 0.5375 59.7275 0.6025 ;
        RECT 61.29 0.445 61.355 0.51 ;
    END
  END rs1_sel[9]
  PIN rs2_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 88.2775 0.69 88.3425 0.825 ;
        RECT 88.0475 0.725 88.3425 0.79 ;
        RECT 88.0475 0.265 88.1125 1.14 ;
    END
  END rs2_rdata
  PIN rs2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.6625 0.505 84.7325 0.64 ;
        RECT 84.5525 0.505 84.7325 0.575 ;
        RECT 84.5525 0.27 84.6225 0.575 ;
        RECT 83.79 0.27 84.6225 0.34 ;
        RECT 83.8825 0.69 83.9525 0.825 ;
        RECT 83.79 0.69 83.9525 0.76 ;
        RECT 83.79 0.27 83.86 0.76 ;
      LAYER metal1 ;
        RECT 84.665 0.505 84.73 0.64 ;
        RECT 83.885 0.69 83.95 0.825 ;
      LAYER via1 ;
        RECT 83.885 0.725 83.95 0.79 ;
        RECT 84.665 0.54 84.73 0.605 ;
    END
  END rs2_sel[0]
  PIN rs2_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 59.105 0.5975 59.245 0.6675 ;
      LAYER metal2 ;
        RECT 58.8475 0.5975 59.245 0.6675 ;
        RECT 58.8475 0.565 58.9175 0.7 ;
      LAYER metal1 ;
        RECT 59.11 0.6 59.245 0.665 ;
        RECT 58.85 0.565 58.915 0.7 ;
      LAYER via2 ;
        RECT 59.14 0.5975 59.21 0.6675 ;
      LAYER via1 ;
        RECT 58.85 0.6 58.915 0.665 ;
        RECT 59.145 0.6 59.21 0.665 ;
    END
  END rs2_sel[10]
  PIN rs2_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 56.405 0.5975 56.545 0.6675 ;
      LAYER metal2 ;
        RECT 56.1475 0.5975 56.545 0.6675 ;
        RECT 56.1475 0.565 56.2175 0.7 ;
      LAYER metal1 ;
        RECT 56.41 0.6 56.545 0.665 ;
        RECT 56.15 0.565 56.215 0.7 ;
      LAYER via2 ;
        RECT 56.44 0.5975 56.51 0.6675 ;
      LAYER via1 ;
        RECT 56.15 0.6 56.215 0.665 ;
        RECT 56.445 0.6 56.51 0.665 ;
    END
  END rs2_sel[11]
  PIN rs2_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 53.705 0.5975 53.845 0.6675 ;
      LAYER metal2 ;
        RECT 53.4475 0.5975 53.845 0.6675 ;
        RECT 53.4475 0.565 53.5175 0.7 ;
      LAYER metal1 ;
        RECT 53.71 0.6 53.845 0.665 ;
        RECT 53.45 0.565 53.515 0.7 ;
      LAYER via2 ;
        RECT 53.74 0.5975 53.81 0.6675 ;
      LAYER via1 ;
        RECT 53.45 0.6 53.515 0.665 ;
        RECT 53.745 0.6 53.81 0.665 ;
    END
  END rs2_sel[12]
  PIN rs2_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 51.005 0.5975 51.145 0.6675 ;
      LAYER metal2 ;
        RECT 50.7475 0.5975 51.145 0.6675 ;
        RECT 50.7475 0.565 50.8175 0.7 ;
      LAYER metal1 ;
        RECT 51.01 0.6 51.145 0.665 ;
        RECT 50.75 0.565 50.815 0.7 ;
      LAYER via2 ;
        RECT 51.04 0.5975 51.11 0.6675 ;
      LAYER via1 ;
        RECT 50.75 0.6 50.815 0.665 ;
        RECT 51.045 0.6 51.11 0.665 ;
    END
  END rs2_sel[13]
  PIN rs2_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 48.305 0.5975 48.445 0.6675 ;
      LAYER metal2 ;
        RECT 48.0475 0.5975 48.445 0.6675 ;
        RECT 48.0475 0.565 48.1175 0.7 ;
      LAYER metal1 ;
        RECT 48.31 0.6 48.445 0.665 ;
        RECT 48.05 0.565 48.115 0.7 ;
      LAYER via2 ;
        RECT 48.34 0.5975 48.41 0.6675 ;
      LAYER via1 ;
        RECT 48.05 0.6 48.115 0.665 ;
        RECT 48.345 0.6 48.41 0.665 ;
    END
  END rs2_sel[14]
  PIN rs2_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 45.605 0.5975 45.745 0.6675 ;
      LAYER metal2 ;
        RECT 45.3475 0.5975 45.745 0.6675 ;
        RECT 45.3475 0.565 45.4175 0.7 ;
      LAYER metal1 ;
        RECT 45.61 0.6 45.745 0.665 ;
        RECT 45.35 0.565 45.415 0.7 ;
      LAYER via2 ;
        RECT 45.64 0.5975 45.71 0.6675 ;
      LAYER via1 ;
        RECT 45.35 0.6 45.415 0.665 ;
        RECT 45.645 0.6 45.71 0.665 ;
    END
  END rs2_sel[15]
  PIN rs2_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 42.905 0.5975 43.045 0.6675 ;
      LAYER metal2 ;
        RECT 42.6475 0.5975 43.045 0.6675 ;
        RECT 42.6475 0.565 42.7175 0.7 ;
      LAYER metal1 ;
        RECT 42.91 0.6 43.045 0.665 ;
        RECT 42.65 0.565 42.715 0.7 ;
      LAYER via2 ;
        RECT 42.94 0.5975 43.01 0.6675 ;
      LAYER via1 ;
        RECT 42.65 0.6 42.715 0.665 ;
        RECT 42.945 0.6 43.01 0.665 ;
    END
  END rs2_sel[16]
  PIN rs2_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 40.205 0.5975 40.345 0.6675 ;
      LAYER metal2 ;
        RECT 39.9475 0.5975 40.345 0.6675 ;
        RECT 39.9475 0.565 40.0175 0.7 ;
      LAYER metal1 ;
        RECT 40.21 0.6 40.345 0.665 ;
        RECT 39.95 0.565 40.015 0.7 ;
      LAYER via2 ;
        RECT 40.24 0.5975 40.31 0.6675 ;
      LAYER via1 ;
        RECT 39.95 0.6 40.015 0.665 ;
        RECT 40.245 0.6 40.31 0.665 ;
    END
  END rs2_sel[17]
  PIN rs2_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 37.505 0.5975 37.645 0.6675 ;
      LAYER metal2 ;
        RECT 37.2475 0.5975 37.645 0.6675 ;
        RECT 37.2475 0.565 37.3175 0.7 ;
      LAYER metal1 ;
        RECT 37.51 0.6 37.645 0.665 ;
        RECT 37.25 0.565 37.315 0.7 ;
      LAYER via2 ;
        RECT 37.54 0.5975 37.61 0.6675 ;
      LAYER via1 ;
        RECT 37.25 0.6 37.315 0.665 ;
        RECT 37.545 0.6 37.61 0.665 ;
    END
  END rs2_sel[18]
  PIN rs2_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 34.805 0.5975 34.945 0.6675 ;
      LAYER metal2 ;
        RECT 34.5475 0.5975 34.945 0.6675 ;
        RECT 34.5475 0.565 34.6175 0.7 ;
      LAYER metal1 ;
        RECT 34.81 0.6 34.945 0.665 ;
        RECT 34.55 0.565 34.615 0.7 ;
      LAYER via2 ;
        RECT 34.84 0.5975 34.91 0.6675 ;
      LAYER via1 ;
        RECT 34.55 0.6 34.615 0.665 ;
        RECT 34.845 0.6 34.91 0.665 ;
    END
  END rs2_sel[19]
  PIN rs2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 83.405 0.5975 83.545 0.6675 ;
      LAYER metal2 ;
        RECT 83.1475 0.5975 83.545 0.6675 ;
        RECT 83.1475 0.565 83.2175 0.7 ;
      LAYER metal1 ;
        RECT 83.41 0.6 83.545 0.665 ;
        RECT 83.15 0.565 83.215 0.7 ;
      LAYER via2 ;
        RECT 83.44 0.5975 83.51 0.6675 ;
      LAYER via1 ;
        RECT 83.15 0.6 83.215 0.665 ;
        RECT 83.445 0.6 83.51 0.665 ;
    END
  END rs2_sel[1]
  PIN rs2_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 32.105 0.5975 32.245 0.6675 ;
      LAYER metal2 ;
        RECT 31.8475 0.5975 32.245 0.6675 ;
        RECT 31.8475 0.565 31.9175 0.7 ;
      LAYER metal1 ;
        RECT 32.11 0.6 32.245 0.665 ;
        RECT 31.85 0.565 31.915 0.7 ;
      LAYER via2 ;
        RECT 32.14 0.5975 32.21 0.6675 ;
      LAYER via1 ;
        RECT 31.85 0.6 31.915 0.665 ;
        RECT 32.145 0.6 32.21 0.665 ;
    END
  END rs2_sel[20]
  PIN rs2_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 29.405 0.5975 29.545 0.6675 ;
      LAYER metal2 ;
        RECT 29.1475 0.5975 29.545 0.6675 ;
        RECT 29.1475 0.565 29.2175 0.7 ;
      LAYER metal1 ;
        RECT 29.41 0.6 29.545 0.665 ;
        RECT 29.15 0.565 29.215 0.7 ;
      LAYER via2 ;
        RECT 29.44 0.5975 29.51 0.6675 ;
      LAYER via1 ;
        RECT 29.15 0.6 29.215 0.665 ;
        RECT 29.445 0.6 29.51 0.665 ;
    END
  END rs2_sel[21]
  PIN rs2_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 26.705 0.5975 26.845 0.6675 ;
      LAYER metal2 ;
        RECT 26.4475 0.5975 26.845 0.6675 ;
        RECT 26.4475 0.565 26.5175 0.7 ;
      LAYER metal1 ;
        RECT 26.71 0.6 26.845 0.665 ;
        RECT 26.45 0.565 26.515 0.7 ;
      LAYER via2 ;
        RECT 26.74 0.5975 26.81 0.6675 ;
      LAYER via1 ;
        RECT 26.45 0.6 26.515 0.665 ;
        RECT 26.745 0.6 26.81 0.665 ;
    END
  END rs2_sel[22]
  PIN rs2_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 24.005 0.5975 24.145 0.6675 ;
      LAYER metal2 ;
        RECT 23.7475 0.5975 24.145 0.6675 ;
        RECT 23.7475 0.565 23.8175 0.7 ;
      LAYER metal1 ;
        RECT 24.01 0.6 24.145 0.665 ;
        RECT 23.75 0.565 23.815 0.7 ;
      LAYER via2 ;
        RECT 24.04 0.5975 24.11 0.6675 ;
      LAYER via1 ;
        RECT 23.75 0.6 23.815 0.665 ;
        RECT 24.045 0.6 24.11 0.665 ;
    END
  END rs2_sel[23]
  PIN rs2_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 21.305 0.5975 21.445 0.6675 ;
      LAYER metal2 ;
        RECT 21.0475 0.5975 21.445 0.6675 ;
        RECT 21.0475 0.565 21.1175 0.7 ;
      LAYER metal1 ;
        RECT 21.31 0.6 21.445 0.665 ;
        RECT 21.05 0.565 21.115 0.7 ;
      LAYER via2 ;
        RECT 21.34 0.5975 21.41 0.6675 ;
      LAYER via1 ;
        RECT 21.05 0.6 21.115 0.665 ;
        RECT 21.345 0.6 21.41 0.665 ;
    END
  END rs2_sel[24]
  PIN rs2_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 18.605 0.5975 18.745 0.6675 ;
      LAYER metal2 ;
        RECT 18.3475 0.5975 18.745 0.6675 ;
        RECT 18.3475 0.565 18.4175 0.7 ;
      LAYER metal1 ;
        RECT 18.61 0.6 18.745 0.665 ;
        RECT 18.35 0.565 18.415 0.7 ;
      LAYER via2 ;
        RECT 18.64 0.5975 18.71 0.6675 ;
      LAYER via1 ;
        RECT 18.35 0.6 18.415 0.665 ;
        RECT 18.645 0.6 18.71 0.665 ;
    END
  END rs2_sel[25]
  PIN rs2_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 15.905 0.5975 16.045 0.6675 ;
      LAYER metal2 ;
        RECT 15.6475 0.5975 16.045 0.6675 ;
        RECT 15.6475 0.565 15.7175 0.7 ;
      LAYER metal1 ;
        RECT 15.91 0.6 16.045 0.665 ;
        RECT 15.65 0.565 15.715 0.7 ;
      LAYER via2 ;
        RECT 15.94 0.5975 16.01 0.6675 ;
      LAYER via1 ;
        RECT 15.65 0.6 15.715 0.665 ;
        RECT 15.945 0.6 16.01 0.665 ;
    END
  END rs2_sel[26]
  PIN rs2_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 13.205 0.5975 13.345 0.6675 ;
      LAYER metal2 ;
        RECT 12.9475 0.5975 13.345 0.6675 ;
        RECT 12.9475 0.565 13.0175 0.7 ;
      LAYER metal1 ;
        RECT 13.21 0.6 13.345 0.665 ;
        RECT 12.95 0.565 13.015 0.7 ;
      LAYER via2 ;
        RECT 13.24 0.5975 13.31 0.6675 ;
      LAYER via1 ;
        RECT 12.95 0.6 13.015 0.665 ;
        RECT 13.245 0.6 13.31 0.665 ;
    END
  END rs2_sel[27]
  PIN rs2_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 10.505 0.5975 10.645 0.6675 ;
      LAYER metal2 ;
        RECT 10.2475 0.5975 10.645 0.6675 ;
        RECT 10.2475 0.565 10.3175 0.7 ;
      LAYER metal1 ;
        RECT 10.51 0.6 10.645 0.665 ;
        RECT 10.25 0.565 10.315 0.7 ;
      LAYER via2 ;
        RECT 10.54 0.5975 10.61 0.6675 ;
      LAYER via1 ;
        RECT 10.25 0.6 10.315 0.665 ;
        RECT 10.545 0.6 10.61 0.665 ;
    END
  END rs2_sel[28]
  PIN rs2_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 7.805 0.5975 7.945 0.6675 ;
      LAYER metal2 ;
        RECT 7.5475 0.5975 7.945 0.6675 ;
        RECT 7.5475 0.565 7.6175 0.7 ;
      LAYER metal1 ;
        RECT 7.81 0.6 7.945 0.665 ;
        RECT 7.55 0.565 7.615 0.7 ;
      LAYER via2 ;
        RECT 7.84 0.5975 7.91 0.6675 ;
      LAYER via1 ;
        RECT 7.55 0.6 7.615 0.665 ;
        RECT 7.845 0.6 7.91 0.665 ;
    END
  END rs2_sel[29]
  PIN rs2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 80.705 0.5975 80.845 0.6675 ;
      LAYER metal2 ;
        RECT 80.4475 0.5975 80.845 0.6675 ;
        RECT 80.4475 0.565 80.5175 0.7 ;
      LAYER metal1 ;
        RECT 80.71 0.6 80.845 0.665 ;
        RECT 80.45 0.565 80.515 0.7 ;
      LAYER via2 ;
        RECT 80.74 0.5975 80.81 0.6675 ;
      LAYER via1 ;
        RECT 80.45 0.6 80.515 0.665 ;
        RECT 80.745 0.6 80.81 0.665 ;
    END
  END rs2_sel[2]
  PIN rs2_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 5.105 0.5975 5.245 0.6675 ;
      LAYER metal2 ;
        RECT 4.8475 0.5975 5.245 0.6675 ;
        RECT 4.8475 0.565 4.9175 0.7 ;
      LAYER metal1 ;
        RECT 5.11 0.6 5.245 0.665 ;
        RECT 4.85 0.565 4.915 0.7 ;
      LAYER via2 ;
        RECT 5.14 0.5975 5.21 0.6675 ;
      LAYER via1 ;
        RECT 4.85 0.6 4.915 0.665 ;
        RECT 5.145 0.6 5.21 0.665 ;
    END
  END rs2_sel[30]
  PIN rs2_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 2.405 0.5975 2.545 0.6675 ;
      LAYER metal2 ;
        RECT 2.1475 0.5975 2.545 0.6675 ;
        RECT 2.1475 0.565 2.2175 0.7 ;
      LAYER metal1 ;
        RECT 2.41 0.6 2.545 0.665 ;
        RECT 2.15 0.565 2.215 0.7 ;
      LAYER via2 ;
        RECT 2.44 0.5975 2.51 0.6675 ;
      LAYER via1 ;
        RECT 2.15 0.6 2.215 0.665 ;
        RECT 2.445 0.6 2.51 0.665 ;
    END
  END rs2_sel[31]
  PIN rs2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 78.005 0.5975 78.145 0.6675 ;
      LAYER metal2 ;
        RECT 77.7475 0.5975 78.145 0.6675 ;
        RECT 77.7475 0.565 77.8175 0.7 ;
      LAYER metal1 ;
        RECT 78.01 0.6 78.145 0.665 ;
        RECT 77.75 0.565 77.815 0.7 ;
      LAYER via2 ;
        RECT 78.04 0.5975 78.11 0.6675 ;
      LAYER via1 ;
        RECT 77.75 0.6 77.815 0.665 ;
        RECT 78.045 0.6 78.11 0.665 ;
    END
  END rs2_sel[3]
  PIN rs2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.305 0.5975 75.445 0.6675 ;
      LAYER metal2 ;
        RECT 75.0475 0.5975 75.445 0.6675 ;
        RECT 75.0475 0.565 75.1175 0.7 ;
      LAYER metal1 ;
        RECT 75.31 0.6 75.445 0.665 ;
        RECT 75.05 0.565 75.115 0.7 ;
      LAYER via2 ;
        RECT 75.34 0.5975 75.41 0.6675 ;
      LAYER via1 ;
        RECT 75.05 0.6 75.115 0.665 ;
        RECT 75.345 0.6 75.41 0.665 ;
    END
  END rs2_sel[4]
  PIN rs2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 72.605 0.5975 72.745 0.6675 ;
      LAYER metal2 ;
        RECT 72.3475 0.5975 72.745 0.6675 ;
        RECT 72.3475 0.565 72.4175 0.7 ;
      LAYER metal1 ;
        RECT 72.61 0.6 72.745 0.665 ;
        RECT 72.35 0.565 72.415 0.7 ;
      LAYER via2 ;
        RECT 72.64 0.5975 72.71 0.6675 ;
      LAYER via1 ;
        RECT 72.35 0.6 72.415 0.665 ;
        RECT 72.645 0.6 72.71 0.665 ;
    END
  END rs2_sel[5]
  PIN rs2_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 69.905 0.5975 70.045 0.6675 ;
      LAYER metal2 ;
        RECT 69.6475 0.5975 70.045 0.6675 ;
        RECT 69.6475 0.565 69.7175 0.7 ;
      LAYER metal1 ;
        RECT 69.91 0.6 70.045 0.665 ;
        RECT 69.65 0.565 69.715 0.7 ;
      LAYER via2 ;
        RECT 69.94 0.5975 70.01 0.6675 ;
      LAYER via1 ;
        RECT 69.65 0.6 69.715 0.665 ;
        RECT 69.945 0.6 70.01 0.665 ;
    END
  END rs2_sel[6]
  PIN rs2_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 67.205 0.5975 67.345 0.6675 ;
      LAYER metal2 ;
        RECT 66.9475 0.5975 67.345 0.6675 ;
        RECT 66.9475 0.565 67.0175 0.7 ;
      LAYER metal1 ;
        RECT 67.21 0.6 67.345 0.665 ;
        RECT 66.95 0.565 67.015 0.7 ;
      LAYER via2 ;
        RECT 67.24 0.5975 67.31 0.6675 ;
      LAYER via1 ;
        RECT 66.95 0.6 67.015 0.665 ;
        RECT 67.245 0.6 67.31 0.665 ;
    END
  END rs2_sel[7]
  PIN rs2_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 64.505 0.5975 64.645 0.6675 ;
      LAYER metal2 ;
        RECT 64.2475 0.5975 64.645 0.6675 ;
        RECT 64.2475 0.565 64.3175 0.7 ;
      LAYER metal1 ;
        RECT 64.51 0.6 64.645 0.665 ;
        RECT 64.25 0.565 64.315 0.7 ;
      LAYER via2 ;
        RECT 64.54 0.5975 64.61 0.6675 ;
      LAYER via1 ;
        RECT 64.25 0.6 64.315 0.665 ;
        RECT 64.545 0.6 64.61 0.665 ;
    END
  END rs2_sel[8]
  PIN rs2_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 61.805 0.5975 61.945 0.6675 ;
      LAYER metal2 ;
        RECT 61.5475 0.5975 61.945 0.6675 ;
        RECT 61.5475 0.565 61.6175 0.7 ;
      LAYER metal1 ;
        RECT 61.81 0.6 61.945 0.665 ;
        RECT 61.55 0.565 61.615 0.7 ;
      LAYER via2 ;
        RECT 61.84 0.5975 61.91 0.6675 ;
      LAYER via1 ;
        RECT 61.55 0.6 61.615 0.665 ;
        RECT 61.845 0.6 61.91 0.665 ;
    END
  END rs2_sel[9]
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.205 88.91 1.405 ;
        RECT 88.235 0.89 88.3 1.405 ;
        RECT 87.4575 0.89 87.5225 1.405 ;
        RECT 87.125 0.89 87.19 1.405 ;
        RECT 86.2375 0.89 86.3025 1.405 ;
        RECT 85.46 0.89 85.525 1.405 ;
        RECT 85.1275 0.89 85.1925 1.405 ;
        RECT 83.9425 0.89 84.0075 1.405 ;
        RECT 83.425 0.89 83.49 1.405 ;
        RECT 82.1675 0.89 82.2325 1.405 ;
        RECT 81.2425 0.89 81.3075 1.405 ;
        RECT 80.725 0.89 80.79 1.405 ;
        RECT 79.4675 0.89 79.5325 1.405 ;
        RECT 78.5425 0.89 78.6075 1.405 ;
        RECT 78.025 0.89 78.09 1.405 ;
        RECT 76.7675 0.89 76.8325 1.405 ;
        RECT 75.8425 0.89 75.9075 1.405 ;
        RECT 75.325 0.89 75.39 1.405 ;
        RECT 74.0675 0.89 74.1325 1.405 ;
        RECT 73.1425 0.89 73.2075 1.405 ;
        RECT 72.625 0.89 72.69 1.405 ;
        RECT 71.3675 0.89 71.4325 1.405 ;
        RECT 70.4425 0.89 70.5075 1.405 ;
        RECT 69.925 0.89 69.99 1.405 ;
        RECT 68.6675 0.89 68.7325 1.405 ;
        RECT 67.7425 0.89 67.8075 1.405 ;
        RECT 67.225 0.89 67.29 1.405 ;
        RECT 65.9675 0.89 66.0325 1.405 ;
        RECT 65.0425 0.89 65.1075 1.405 ;
        RECT 64.525 0.89 64.59 1.405 ;
        RECT 63.2675 0.89 63.3325 1.405 ;
        RECT 62.3425 0.89 62.4075 1.405 ;
        RECT 61.825 0.89 61.89 1.405 ;
        RECT 60.5675 0.89 60.6325 1.405 ;
        RECT 59.6425 0.89 59.7075 1.405 ;
        RECT 59.125 0.89 59.19 1.405 ;
        RECT 57.8675 0.89 57.9325 1.405 ;
        RECT 56.9425 0.89 57.0075 1.405 ;
        RECT 56.425 0.89 56.49 1.405 ;
        RECT 55.1675 0.89 55.2325 1.405 ;
        RECT 54.2425 0.89 54.3075 1.405 ;
        RECT 53.725 0.89 53.79 1.405 ;
        RECT 52.4675 0.89 52.5325 1.405 ;
        RECT 51.5425 0.89 51.6075 1.405 ;
        RECT 51.025 0.89 51.09 1.405 ;
        RECT 49.7675 0.89 49.8325 1.405 ;
        RECT 48.8425 0.89 48.9075 1.405 ;
        RECT 48.325 0.89 48.39 1.405 ;
        RECT 47.0675 0.89 47.1325 1.405 ;
        RECT 46.1425 0.89 46.2075 1.405 ;
        RECT 45.625 0.89 45.69 1.405 ;
        RECT 44.3675 0.89 44.4325 1.405 ;
        RECT 43.4425 0.89 43.5075 1.405 ;
        RECT 42.925 0.89 42.99 1.405 ;
        RECT 41.6675 0.89 41.7325 1.405 ;
        RECT 40.7425 0.89 40.8075 1.405 ;
        RECT 40.225 0.89 40.29 1.405 ;
        RECT 38.9675 0.89 39.0325 1.405 ;
        RECT 38.0425 0.89 38.1075 1.405 ;
        RECT 37.525 0.89 37.59 1.405 ;
        RECT 36.2675 0.89 36.3325 1.405 ;
        RECT 35.3425 0.89 35.4075 1.405 ;
        RECT 34.825 0.89 34.89 1.405 ;
        RECT 33.5675 0.89 33.6325 1.405 ;
        RECT 32.6425 0.89 32.7075 1.405 ;
        RECT 32.125 0.89 32.19 1.405 ;
        RECT 30.8675 0.89 30.9325 1.405 ;
        RECT 29.9425 0.89 30.0075 1.405 ;
        RECT 29.425 0.89 29.49 1.405 ;
        RECT 28.1675 0.89 28.2325 1.405 ;
        RECT 27.2425 0.89 27.3075 1.405 ;
        RECT 26.725 0.89 26.79 1.405 ;
        RECT 25.4675 0.89 25.5325 1.405 ;
        RECT 24.5425 0.89 24.6075 1.405 ;
        RECT 24.025 0.89 24.09 1.405 ;
        RECT 22.7675 0.89 22.8325 1.405 ;
        RECT 21.8425 0.89 21.9075 1.405 ;
        RECT 21.325 0.89 21.39 1.405 ;
        RECT 20.0675 0.89 20.1325 1.405 ;
        RECT 19.1425 0.89 19.2075 1.405 ;
        RECT 18.625 0.89 18.69 1.405 ;
        RECT 17.3675 0.89 17.4325 1.405 ;
        RECT 16.4425 0.89 16.5075 1.405 ;
        RECT 15.925 0.89 15.99 1.405 ;
        RECT 14.6675 0.89 14.7325 1.405 ;
        RECT 13.7425 0.89 13.8075 1.405 ;
        RECT 13.225 0.89 13.29 1.405 ;
        RECT 11.9675 0.89 12.0325 1.405 ;
        RECT 11.0425 0.89 11.1075 1.405 ;
        RECT 10.525 0.89 10.59 1.405 ;
        RECT 9.2675 0.89 9.3325 1.405 ;
        RECT 8.3425 0.89 8.4075 1.405 ;
        RECT 7.825 0.89 7.89 1.405 ;
        RECT 6.5675 0.89 6.6325 1.405 ;
        RECT 5.6425 0.89 5.7075 1.405 ;
        RECT 5.125 0.89 5.19 1.405 ;
        RECT 3.8675 0.89 3.9325 1.405 ;
        RECT 2.9425 0.89 3.0075 1.405 ;
        RECT 2.425 0.89 2.49 1.405 ;
        RECT 1.1675 0.89 1.2325 1.405 ;
        RECT 0.2425 0.89 0.3075 1.405 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 88.91 0.2 ;
        RECT 88.2325 0 88.2975 0.425 ;
        RECT 87.4575 0 87.5225 0.425 ;
        RECT 87.125 0 87.19 0.425 ;
        RECT 86.235 0 86.3 0.425 ;
        RECT 85.46 0 85.525 0.425 ;
        RECT 85.1275 0 85.1925 0.425 ;
        RECT 84.535 0 84.6 1.14 ;
        RECT 83.9425 0 84.0075 0.425 ;
        RECT 83.425 0 83.49 0.425 ;
        RECT 82.1675 0 82.2325 0.425 ;
        RECT 81.2425 0 81.3075 0.425 ;
        RECT 80.725 0 80.79 0.425 ;
        RECT 79.4675 0 79.5325 0.425 ;
        RECT 78.5425 0 78.6075 0.425 ;
        RECT 78.025 0 78.09 0.425 ;
        RECT 76.7675 0 76.8325 0.425 ;
        RECT 75.8425 0 75.9075 0.425 ;
        RECT 75.325 0 75.39 0.425 ;
        RECT 74.0675 0 74.1325 0.425 ;
        RECT 73.1425 0 73.2075 0.425 ;
        RECT 72.625 0 72.69 0.425 ;
        RECT 71.3675 0 71.4325 0.425 ;
        RECT 70.4425 0 70.5075 0.425 ;
        RECT 69.925 0 69.99 0.425 ;
        RECT 68.6675 0 68.7325 0.425 ;
        RECT 67.7425 0 67.8075 0.425 ;
        RECT 67.225 0 67.29 0.425 ;
        RECT 65.9675 0 66.0325 0.425 ;
        RECT 65.0425 0 65.1075 0.425 ;
        RECT 64.525 0 64.59 0.425 ;
        RECT 63.2675 0 63.3325 0.425 ;
        RECT 62.3425 0 62.4075 0.425 ;
        RECT 61.825 0 61.89 0.425 ;
        RECT 60.5675 0 60.6325 0.425 ;
        RECT 59.6425 0 59.7075 0.425 ;
        RECT 59.125 0 59.19 0.425 ;
        RECT 57.8675 0 57.9325 0.425 ;
        RECT 56.9425 0 57.0075 0.425 ;
        RECT 56.425 0 56.49 0.425 ;
        RECT 55.1675 0 55.2325 0.425 ;
        RECT 54.2425 0 54.3075 0.425 ;
        RECT 53.725 0 53.79 0.425 ;
        RECT 52.4675 0 52.5325 0.425 ;
        RECT 51.5425 0 51.6075 0.425 ;
        RECT 51.025 0 51.09 0.425 ;
        RECT 49.7675 0 49.8325 0.425 ;
        RECT 48.8425 0 48.9075 0.425 ;
        RECT 48.325 0 48.39 0.425 ;
        RECT 47.0675 0 47.1325 0.425 ;
        RECT 46.1425 0 46.2075 0.425 ;
        RECT 45.625 0 45.69 0.425 ;
        RECT 44.3675 0 44.4325 0.425 ;
        RECT 43.4425 0 43.5075 0.425 ;
        RECT 42.925 0 42.99 0.425 ;
        RECT 41.6675 0 41.7325 0.425 ;
        RECT 40.7425 0 40.8075 0.425 ;
        RECT 40.225 0 40.29 0.425 ;
        RECT 38.9675 0 39.0325 0.425 ;
        RECT 38.0425 0 38.1075 0.425 ;
        RECT 37.525 0 37.59 0.425 ;
        RECT 36.2675 0 36.3325 0.425 ;
        RECT 35.3425 0 35.4075 0.425 ;
        RECT 34.825 0 34.89 0.425 ;
        RECT 33.5675 0 33.6325 0.425 ;
        RECT 32.6425 0 32.7075 0.425 ;
        RECT 32.125 0 32.19 0.425 ;
        RECT 30.8675 0 30.9325 0.425 ;
        RECT 29.9425 0 30.0075 0.425 ;
        RECT 29.425 0 29.49 0.425 ;
        RECT 28.1675 0 28.2325 0.425 ;
        RECT 27.2425 0 27.3075 0.425 ;
        RECT 26.725 0 26.79 0.425 ;
        RECT 25.4675 0 25.5325 0.425 ;
        RECT 24.5425 0 24.6075 0.425 ;
        RECT 24.025 0 24.09 0.425 ;
        RECT 22.7675 0 22.8325 0.425 ;
        RECT 21.8425 0 21.9075 0.425 ;
        RECT 21.325 0 21.39 0.425 ;
        RECT 20.0675 0 20.1325 0.425 ;
        RECT 19.1425 0 19.2075 0.425 ;
        RECT 18.625 0 18.69 0.425 ;
        RECT 17.3675 0 17.4325 0.425 ;
        RECT 16.4425 0 16.5075 0.425 ;
        RECT 15.925 0 15.99 0.425 ;
        RECT 14.6675 0 14.7325 0.425 ;
        RECT 13.7425 0 13.8075 0.425 ;
        RECT 13.225 0 13.29 0.425 ;
        RECT 11.9675 0 12.0325 0.425 ;
        RECT 11.0425 0 11.1075 0.425 ;
        RECT 10.525 0 10.59 0.425 ;
        RECT 9.2675 0 9.3325 0.425 ;
        RECT 8.3425 0 8.4075 0.425 ;
        RECT 7.825 0 7.89 0.425 ;
        RECT 6.5675 0 6.6325 0.425 ;
        RECT 5.6425 0 5.7075 0.425 ;
        RECT 5.125 0 5.19 0.425 ;
        RECT 3.8675 0 3.9325 0.425 ;
        RECT 2.9425 0 3.0075 0.425 ;
        RECT 2.425 0 2.49 0.425 ;
        RECT 1.1675 0 1.2325 0.425 ;
        RECT 0.2425 0 0.3075 0.425 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 88.79 0.265 88.855 1.14 ;
      RECT 88.79 0.5825 88.8625 0.7175 ;
      RECT 88.1925 0.56 88.3275 0.625 ;
      RECT 88.1925 0.49 88.2575 0.625 ;
      RECT 87.9025 0.265 87.9675 1.14 ;
      RECT 87.9025 0.5825 87.9775 0.7175 ;
      RECT 87.3125 0.265 87.3775 1.14 ;
      RECT 87.0675 0.49 87.1325 0.625 ;
      RECT 87.0675 0.525 87.3775 0.59 ;
      RECT 86.7925 0.265 86.8575 1.14 ;
      RECT 86.7925 0.5825 86.865 0.7175 ;
      RECT 86.195 0.56 86.33 0.625 ;
      RECT 86.195 0.49 86.26 0.625 ;
      RECT 85.905 0.265 85.97 1.14 ;
      RECT 85.905 0.5825 85.98 0.7175 ;
      RECT 85.315 0.265 85.38 1.14 ;
      RECT 85.07 0.49 85.135 0.625 ;
      RECT 85.07 0.525 85.38 0.59 ;
      RECT 84.795 0.265 84.86 1.14 ;
      RECT 84.725 0.265 84.86 0.33 ;
      RECT 84.275 0.265 84.34 1.14 ;
      RECT 84.275 0.625 84.4675 0.69 ;
      RECT 83.28 0.265 83.345 1.14 ;
      RECT 83.21 0.265 83.345 0.33 ;
      RECT 83.02 0.265 83.085 1.14 ;
      RECT 82.9475 0.265 83.085 0.33 ;
      RECT 82.76 0.265 82.825 1.14 ;
      RECT 82.76 0.625 82.955 0.69 ;
      RECT 82.615 0.265 82.68 1.14 ;
      RECT 82.485 0.9775 82.68 1.0425 ;
      RECT 82.355 0.265 82.42 1.14 ;
      RECT 82.355 0.265 82.49 0.33 ;
      RECT 81.98 0.265 82.045 1.14 ;
      RECT 82.22 0.49 82.285 0.625 ;
      RECT 81.98 0.525 82.285 0.59 ;
      RECT 81.835 0.265 81.9 1.14 ;
      RECT 81.765 0.9775 81.9 1.0425 ;
      RECT 80.58 0.265 80.645 1.14 ;
      RECT 80.51 0.265 80.645 0.33 ;
      RECT 80.32 0.265 80.385 1.14 ;
      RECT 80.2475 0.265 80.385 0.33 ;
      RECT 80.06 0.265 80.125 1.14 ;
      RECT 80.06 0.625 80.255 0.69 ;
      RECT 79.915 0.265 79.98 1.14 ;
      RECT 79.785 0.9775 79.98 1.0425 ;
      RECT 79.655 0.265 79.72 1.14 ;
      RECT 79.655 0.265 79.79 0.33 ;
      RECT 79.28 0.265 79.345 1.14 ;
      RECT 79.52 0.49 79.585 0.625 ;
      RECT 79.28 0.525 79.585 0.59 ;
      RECT 79.135 0.265 79.2 1.14 ;
      RECT 79.065 0.9775 79.2 1.0425 ;
      RECT 77.88 0.265 77.945 1.14 ;
      RECT 77.81 0.265 77.945 0.33 ;
      RECT 77.62 0.265 77.685 1.14 ;
      RECT 77.5475 0.265 77.685 0.33 ;
      RECT 77.36 0.265 77.425 1.14 ;
      RECT 77.36 0.625 77.555 0.69 ;
      RECT 77.215 0.265 77.28 1.14 ;
      RECT 77.085 0.9775 77.28 1.0425 ;
      RECT 76.955 0.265 77.02 1.14 ;
      RECT 76.955 0.265 77.09 0.33 ;
      RECT 76.58 0.265 76.645 1.14 ;
      RECT 76.82 0.49 76.885 0.625 ;
      RECT 76.58 0.525 76.885 0.59 ;
      RECT 76.435 0.265 76.5 1.14 ;
      RECT 76.365 0.9775 76.5 1.0425 ;
      RECT 75.18 0.265 75.245 1.14 ;
      RECT 75.11 0.265 75.245 0.33 ;
      RECT 74.92 0.265 74.985 1.14 ;
      RECT 74.8475 0.265 74.985 0.33 ;
      RECT 74.66 0.265 74.725 1.14 ;
      RECT 74.66 0.625 74.855 0.69 ;
      RECT 74.515 0.265 74.58 1.14 ;
      RECT 74.385 0.9775 74.58 1.0425 ;
      RECT 74.255 0.265 74.32 1.14 ;
      RECT 74.255 0.265 74.39 0.33 ;
      RECT 73.88 0.265 73.945 1.14 ;
      RECT 74.12 0.49 74.185 0.625 ;
      RECT 73.88 0.525 74.185 0.59 ;
      RECT 73.735 0.265 73.8 1.14 ;
      RECT 73.665 0.9775 73.8 1.0425 ;
      RECT 72.48 0.265 72.545 1.14 ;
      RECT 72.41 0.265 72.545 0.33 ;
      RECT 72.22 0.265 72.285 1.14 ;
      RECT 72.1475 0.265 72.285 0.33 ;
      RECT 71.96 0.265 72.025 1.14 ;
      RECT 71.96 0.625 72.155 0.69 ;
      RECT 71.815 0.265 71.88 1.14 ;
      RECT 71.685 0.9775 71.88 1.0425 ;
      RECT 71.555 0.265 71.62 1.14 ;
      RECT 71.555 0.265 71.69 0.33 ;
      RECT 71.18 0.265 71.245 1.14 ;
      RECT 71.42 0.49 71.485 0.625 ;
      RECT 71.18 0.525 71.485 0.59 ;
      RECT 71.035 0.265 71.1 1.14 ;
      RECT 70.965 0.9775 71.1 1.0425 ;
      RECT 69.78 0.265 69.845 1.14 ;
      RECT 69.71 0.265 69.845 0.33 ;
      RECT 69.52 0.265 69.585 1.14 ;
      RECT 69.4475 0.265 69.585 0.33 ;
      RECT 69.26 0.265 69.325 1.14 ;
      RECT 69.26 0.625 69.455 0.69 ;
      RECT 69.115 0.265 69.18 1.14 ;
      RECT 68.985 0.9775 69.18 1.0425 ;
      RECT 68.855 0.265 68.92 1.14 ;
      RECT 68.855 0.265 68.99 0.33 ;
      RECT 68.48 0.265 68.545 1.14 ;
      RECT 68.72 0.49 68.785 0.625 ;
      RECT 68.48 0.525 68.785 0.59 ;
      RECT 68.335 0.265 68.4 1.14 ;
      RECT 68.265 0.9775 68.4 1.0425 ;
      RECT 67.08 0.265 67.145 1.14 ;
      RECT 67.01 0.265 67.145 0.33 ;
      RECT 66.82 0.265 66.885 1.14 ;
      RECT 66.7475 0.265 66.885 0.33 ;
      RECT 66.56 0.265 66.625 1.14 ;
      RECT 66.56 0.625 66.755 0.69 ;
      RECT 66.415 0.265 66.48 1.14 ;
      RECT 66.285 0.9775 66.48 1.0425 ;
      RECT 66.155 0.265 66.22 1.14 ;
      RECT 66.155 0.265 66.29 0.33 ;
      RECT 65.78 0.265 65.845 1.14 ;
      RECT 66.02 0.49 66.085 0.625 ;
      RECT 65.78 0.525 66.085 0.59 ;
      RECT 65.635 0.265 65.7 1.14 ;
      RECT 65.565 0.9775 65.7 1.0425 ;
      RECT 64.38 0.265 64.445 1.14 ;
      RECT 64.31 0.265 64.445 0.33 ;
      RECT 64.12 0.265 64.185 1.14 ;
      RECT 64.0475 0.265 64.185 0.33 ;
      RECT 63.86 0.265 63.925 1.14 ;
      RECT 63.86 0.625 64.055 0.69 ;
      RECT 63.715 0.265 63.78 1.14 ;
      RECT 63.585 0.9775 63.78 1.0425 ;
      RECT 63.455 0.265 63.52 1.14 ;
      RECT 63.455 0.265 63.59 0.33 ;
      RECT 63.08 0.265 63.145 1.14 ;
      RECT 63.32 0.49 63.385 0.625 ;
      RECT 63.08 0.525 63.385 0.59 ;
      RECT 62.935 0.265 63 1.14 ;
      RECT 62.865 0.9775 63 1.0425 ;
      RECT 61.68 0.265 61.745 1.14 ;
      RECT 61.61 0.265 61.745 0.33 ;
      RECT 61.42 0.265 61.485 1.14 ;
      RECT 61.3475 0.265 61.485 0.33 ;
      RECT 61.16 0.265 61.225 1.14 ;
      RECT 61.16 0.625 61.355 0.69 ;
      RECT 61.015 0.265 61.08 1.14 ;
      RECT 60.885 0.9775 61.08 1.0425 ;
      RECT 60.755 0.265 60.82 1.14 ;
      RECT 60.755 0.265 60.89 0.33 ;
      RECT 60.38 0.265 60.445 1.14 ;
      RECT 60.62 0.49 60.685 0.625 ;
      RECT 60.38 0.525 60.685 0.59 ;
      RECT 60.235 0.265 60.3 1.14 ;
      RECT 60.165 0.9775 60.3 1.0425 ;
      RECT 58.98 0.265 59.045 1.14 ;
      RECT 58.91 0.265 59.045 0.33 ;
      RECT 58.72 0.265 58.785 1.14 ;
      RECT 58.6475 0.265 58.785 0.33 ;
      RECT 58.46 0.265 58.525 1.14 ;
      RECT 58.46 0.625 58.655 0.69 ;
      RECT 58.315 0.265 58.38 1.14 ;
      RECT 58.185 0.9775 58.38 1.0425 ;
      RECT 58.055 0.265 58.12 1.14 ;
      RECT 58.055 0.265 58.19 0.33 ;
      RECT 57.68 0.265 57.745 1.14 ;
      RECT 57.92 0.49 57.985 0.625 ;
      RECT 57.68 0.525 57.985 0.59 ;
      RECT 57.535 0.265 57.6 1.14 ;
      RECT 57.465 0.9775 57.6 1.0425 ;
      RECT 56.28 0.265 56.345 1.14 ;
      RECT 56.21 0.265 56.345 0.33 ;
      RECT 56.02 0.265 56.085 1.14 ;
      RECT 55.9475 0.265 56.085 0.33 ;
      RECT 55.76 0.265 55.825 1.14 ;
      RECT 55.76 0.625 55.955 0.69 ;
      RECT 55.615 0.265 55.68 1.14 ;
      RECT 55.485 0.9775 55.68 1.0425 ;
      RECT 55.355 0.265 55.42 1.14 ;
      RECT 55.355 0.265 55.49 0.33 ;
      RECT 54.98 0.265 55.045 1.14 ;
      RECT 55.22 0.49 55.285 0.625 ;
      RECT 54.98 0.525 55.285 0.59 ;
      RECT 54.835 0.265 54.9 1.14 ;
      RECT 54.765 0.9775 54.9 1.0425 ;
      RECT 53.58 0.265 53.645 1.14 ;
      RECT 53.51 0.265 53.645 0.33 ;
      RECT 53.32 0.265 53.385 1.14 ;
      RECT 53.2475 0.265 53.385 0.33 ;
      RECT 53.06 0.265 53.125 1.14 ;
      RECT 53.06 0.625 53.255 0.69 ;
      RECT 52.915 0.265 52.98 1.14 ;
      RECT 52.785 0.9775 52.98 1.0425 ;
      RECT 52.655 0.265 52.72 1.14 ;
      RECT 52.655 0.265 52.79 0.33 ;
      RECT 52.28 0.265 52.345 1.14 ;
      RECT 52.52 0.49 52.585 0.625 ;
      RECT 52.28 0.525 52.585 0.59 ;
      RECT 52.135 0.265 52.2 1.14 ;
      RECT 52.065 0.9775 52.2 1.0425 ;
      RECT 50.88 0.265 50.945 1.14 ;
      RECT 50.81 0.265 50.945 0.33 ;
      RECT 50.62 0.265 50.685 1.14 ;
      RECT 50.5475 0.265 50.685 0.33 ;
      RECT 50.36 0.265 50.425 1.14 ;
      RECT 50.36 0.625 50.555 0.69 ;
      RECT 50.215 0.265 50.28 1.14 ;
      RECT 50.085 0.9775 50.28 1.0425 ;
      RECT 49.955 0.265 50.02 1.14 ;
      RECT 49.955 0.265 50.09 0.33 ;
      RECT 49.58 0.265 49.645 1.14 ;
      RECT 49.82 0.49 49.885 0.625 ;
      RECT 49.58 0.525 49.885 0.59 ;
      RECT 49.435 0.265 49.5 1.14 ;
      RECT 49.365 0.9775 49.5 1.0425 ;
      RECT 48.18 0.265 48.245 1.14 ;
      RECT 48.11 0.265 48.245 0.33 ;
      RECT 47.92 0.265 47.985 1.14 ;
      RECT 47.8475 0.265 47.985 0.33 ;
      RECT 47.66 0.265 47.725 1.14 ;
      RECT 47.66 0.625 47.855 0.69 ;
      RECT 47.515 0.265 47.58 1.14 ;
      RECT 47.385 0.9775 47.58 1.0425 ;
      RECT 47.255 0.265 47.32 1.14 ;
      RECT 47.255 0.265 47.39 0.33 ;
      RECT 46.88 0.265 46.945 1.14 ;
      RECT 47.12 0.49 47.185 0.625 ;
      RECT 46.88 0.525 47.185 0.59 ;
      RECT 46.735 0.265 46.8 1.14 ;
      RECT 46.665 0.9775 46.8 1.0425 ;
      RECT 45.48 0.265 45.545 1.14 ;
      RECT 45.41 0.265 45.545 0.33 ;
      RECT 45.22 0.265 45.285 1.14 ;
      RECT 45.1475 0.265 45.285 0.33 ;
      RECT 44.96 0.265 45.025 1.14 ;
      RECT 44.96 0.625 45.155 0.69 ;
      RECT 44.815 0.265 44.88 1.14 ;
      RECT 44.685 0.9775 44.88 1.0425 ;
      RECT 44.555 0.265 44.62 1.14 ;
      RECT 44.555 0.265 44.69 0.33 ;
      RECT 44.18 0.265 44.245 1.14 ;
      RECT 44.42 0.49 44.485 0.625 ;
      RECT 44.18 0.525 44.485 0.59 ;
      RECT 44.035 0.265 44.1 1.14 ;
      RECT 43.965 0.9775 44.1 1.0425 ;
      RECT 42.78 0.265 42.845 1.14 ;
      RECT 42.71 0.265 42.845 0.33 ;
      RECT 42.52 0.265 42.585 1.14 ;
      RECT 42.4475 0.265 42.585 0.33 ;
      RECT 42.26 0.265 42.325 1.14 ;
      RECT 42.26 0.625 42.455 0.69 ;
      RECT 42.115 0.265 42.18 1.14 ;
      RECT 41.985 0.9775 42.18 1.0425 ;
      RECT 41.855 0.265 41.92 1.14 ;
      RECT 41.855 0.265 41.99 0.33 ;
      RECT 41.48 0.265 41.545 1.14 ;
      RECT 41.72 0.49 41.785 0.625 ;
      RECT 41.48 0.525 41.785 0.59 ;
      RECT 41.335 0.265 41.4 1.14 ;
      RECT 41.265 0.9775 41.4 1.0425 ;
      RECT 40.08 0.265 40.145 1.14 ;
      RECT 40.01 0.265 40.145 0.33 ;
      RECT 39.82 0.265 39.885 1.14 ;
      RECT 39.7475 0.265 39.885 0.33 ;
      RECT 39.56 0.265 39.625 1.14 ;
      RECT 39.56 0.625 39.755 0.69 ;
      RECT 39.415 0.265 39.48 1.14 ;
      RECT 39.285 0.9775 39.48 1.0425 ;
      RECT 39.155 0.265 39.22 1.14 ;
      RECT 39.155 0.265 39.29 0.33 ;
      RECT 38.78 0.265 38.845 1.14 ;
      RECT 39.02 0.49 39.085 0.625 ;
      RECT 38.78 0.525 39.085 0.59 ;
      RECT 38.635 0.265 38.7 1.14 ;
      RECT 38.565 0.9775 38.7 1.0425 ;
      RECT 37.38 0.265 37.445 1.14 ;
      RECT 37.31 0.265 37.445 0.33 ;
      RECT 37.12 0.265 37.185 1.14 ;
      RECT 37.0475 0.265 37.185 0.33 ;
      RECT 36.86 0.265 36.925 1.14 ;
      RECT 36.86 0.625 37.055 0.69 ;
      RECT 36.715 0.265 36.78 1.14 ;
      RECT 36.585 0.9775 36.78 1.0425 ;
      RECT 36.455 0.265 36.52 1.14 ;
      RECT 36.455 0.265 36.59 0.33 ;
      RECT 36.08 0.265 36.145 1.14 ;
      RECT 36.32 0.49 36.385 0.625 ;
      RECT 36.08 0.525 36.385 0.59 ;
      RECT 35.935 0.265 36 1.14 ;
      RECT 35.865 0.9775 36 1.0425 ;
      RECT 34.68 0.265 34.745 1.14 ;
      RECT 34.61 0.265 34.745 0.33 ;
      RECT 34.42 0.265 34.485 1.14 ;
      RECT 34.3475 0.265 34.485 0.33 ;
      RECT 34.16 0.265 34.225 1.14 ;
      RECT 34.16 0.625 34.355 0.69 ;
      RECT 34.015 0.265 34.08 1.14 ;
      RECT 33.885 0.9775 34.08 1.0425 ;
      RECT 33.755 0.265 33.82 1.14 ;
      RECT 33.755 0.265 33.89 0.33 ;
      RECT 33.38 0.265 33.445 1.14 ;
      RECT 33.62 0.49 33.685 0.625 ;
      RECT 33.38 0.525 33.685 0.59 ;
      RECT 33.235 0.265 33.3 1.14 ;
      RECT 33.165 0.9775 33.3 1.0425 ;
      RECT 31.98 0.265 32.045 1.14 ;
      RECT 31.91 0.265 32.045 0.33 ;
      RECT 31.72 0.265 31.785 1.14 ;
      RECT 31.6475 0.265 31.785 0.33 ;
      RECT 31.46 0.265 31.525 1.14 ;
      RECT 31.46 0.625 31.655 0.69 ;
      RECT 31.315 0.265 31.38 1.14 ;
      RECT 31.185 0.9775 31.38 1.0425 ;
      RECT 31.055 0.265 31.12 1.14 ;
      RECT 31.055 0.265 31.19 0.33 ;
      RECT 30.68 0.265 30.745 1.14 ;
      RECT 30.92 0.49 30.985 0.625 ;
      RECT 30.68 0.525 30.985 0.59 ;
      RECT 30.535 0.265 30.6 1.14 ;
      RECT 30.465 0.9775 30.6 1.0425 ;
      RECT 29.28 0.265 29.345 1.14 ;
      RECT 29.21 0.265 29.345 0.33 ;
      RECT 29.02 0.265 29.085 1.14 ;
      RECT 28.9475 0.265 29.085 0.33 ;
      RECT 28.76 0.265 28.825 1.14 ;
      RECT 28.76 0.625 28.955 0.69 ;
      RECT 28.615 0.265 28.68 1.14 ;
      RECT 28.485 0.9775 28.68 1.0425 ;
      RECT 28.355 0.265 28.42 1.14 ;
      RECT 28.355 0.265 28.49 0.33 ;
      RECT 27.98 0.265 28.045 1.14 ;
      RECT 28.22 0.49 28.285 0.625 ;
      RECT 27.98 0.525 28.285 0.59 ;
      RECT 27.835 0.265 27.9 1.14 ;
      RECT 27.765 0.9775 27.9 1.0425 ;
      RECT 26.58 0.265 26.645 1.14 ;
      RECT 26.51 0.265 26.645 0.33 ;
      RECT 26.32 0.265 26.385 1.14 ;
      RECT 26.2475 0.265 26.385 0.33 ;
      RECT 26.06 0.265 26.125 1.14 ;
      RECT 26.06 0.625 26.255 0.69 ;
      RECT 25.915 0.265 25.98 1.14 ;
      RECT 25.785 0.9775 25.98 1.0425 ;
      RECT 25.655 0.265 25.72 1.14 ;
      RECT 25.655 0.265 25.79 0.33 ;
      RECT 25.28 0.265 25.345 1.14 ;
      RECT 25.52 0.49 25.585 0.625 ;
      RECT 25.28 0.525 25.585 0.59 ;
      RECT 25.135 0.265 25.2 1.14 ;
      RECT 25.065 0.9775 25.2 1.0425 ;
      RECT 23.88 0.265 23.945 1.14 ;
      RECT 23.81 0.265 23.945 0.33 ;
      RECT 23.62 0.265 23.685 1.14 ;
      RECT 23.5475 0.265 23.685 0.33 ;
      RECT 23.36 0.265 23.425 1.14 ;
      RECT 23.36 0.625 23.555 0.69 ;
      RECT 23.215 0.265 23.28 1.14 ;
      RECT 23.085 0.9775 23.28 1.0425 ;
      RECT 22.955 0.265 23.02 1.14 ;
      RECT 22.955 0.265 23.09 0.33 ;
      RECT 22.58 0.265 22.645 1.14 ;
      RECT 22.82 0.49 22.885 0.625 ;
      RECT 22.58 0.525 22.885 0.59 ;
      RECT 22.435 0.265 22.5 1.14 ;
      RECT 22.365 0.9775 22.5 1.0425 ;
      RECT 21.18 0.265 21.245 1.14 ;
      RECT 21.11 0.265 21.245 0.33 ;
      RECT 20.92 0.265 20.985 1.14 ;
      RECT 20.8475 0.265 20.985 0.33 ;
      RECT 20.66 0.265 20.725 1.14 ;
      RECT 20.66 0.625 20.855 0.69 ;
      RECT 20.515 0.265 20.58 1.14 ;
      RECT 20.385 0.9775 20.58 1.0425 ;
      RECT 20.255 0.265 20.32 1.14 ;
      RECT 20.255 0.265 20.39 0.33 ;
      RECT 19.88 0.265 19.945 1.14 ;
      RECT 20.12 0.49 20.185 0.625 ;
      RECT 19.88 0.525 20.185 0.59 ;
      RECT 19.735 0.265 19.8 1.14 ;
      RECT 19.665 0.9775 19.8 1.0425 ;
      RECT 18.48 0.265 18.545 1.14 ;
      RECT 18.41 0.265 18.545 0.33 ;
      RECT 18.22 0.265 18.285 1.14 ;
      RECT 18.1475 0.265 18.285 0.33 ;
      RECT 17.96 0.265 18.025 1.14 ;
      RECT 17.96 0.625 18.155 0.69 ;
      RECT 17.815 0.265 17.88 1.14 ;
      RECT 17.685 0.9775 17.88 1.0425 ;
      RECT 17.555 0.265 17.62 1.14 ;
      RECT 17.555 0.265 17.69 0.33 ;
      RECT 17.18 0.265 17.245 1.14 ;
      RECT 17.42 0.49 17.485 0.625 ;
      RECT 17.18 0.525 17.485 0.59 ;
      RECT 17.035 0.265 17.1 1.14 ;
      RECT 16.965 0.9775 17.1 1.0425 ;
      RECT 15.78 0.265 15.845 1.14 ;
      RECT 15.71 0.265 15.845 0.33 ;
      RECT 15.52 0.265 15.585 1.14 ;
      RECT 15.4475 0.265 15.585 0.33 ;
      RECT 15.26 0.265 15.325 1.14 ;
      RECT 15.26 0.625 15.455 0.69 ;
      RECT 15.115 0.265 15.18 1.14 ;
      RECT 14.985 0.9775 15.18 1.0425 ;
      RECT 14.855 0.265 14.92 1.14 ;
      RECT 14.855 0.265 14.99 0.33 ;
      RECT 14.48 0.265 14.545 1.14 ;
      RECT 14.72 0.49 14.785 0.625 ;
      RECT 14.48 0.525 14.785 0.59 ;
      RECT 14.335 0.265 14.4 1.14 ;
      RECT 14.265 0.9775 14.4 1.0425 ;
      RECT 13.08 0.265 13.145 1.14 ;
      RECT 13.01 0.265 13.145 0.33 ;
      RECT 12.82 0.265 12.885 1.14 ;
      RECT 12.7475 0.265 12.885 0.33 ;
      RECT 12.56 0.265 12.625 1.14 ;
      RECT 12.56 0.625 12.755 0.69 ;
      RECT 12.415 0.265 12.48 1.14 ;
      RECT 12.285 0.9775 12.48 1.0425 ;
      RECT 12.155 0.265 12.22 1.14 ;
      RECT 12.155 0.265 12.29 0.33 ;
      RECT 11.78 0.265 11.845 1.14 ;
      RECT 12.02 0.49 12.085 0.625 ;
      RECT 11.78 0.525 12.085 0.59 ;
      RECT 11.635 0.265 11.7 1.14 ;
      RECT 11.565 0.9775 11.7 1.0425 ;
      RECT 10.38 0.265 10.445 1.14 ;
      RECT 10.31 0.265 10.445 0.33 ;
      RECT 10.12 0.265 10.185 1.14 ;
      RECT 10.0475 0.265 10.185 0.33 ;
      RECT 9.86 0.265 9.925 1.14 ;
      RECT 9.86 0.625 10.055 0.69 ;
      RECT 9.715 0.265 9.78 1.14 ;
      RECT 9.585 0.9775 9.78 1.0425 ;
      RECT 9.455 0.265 9.52 1.14 ;
      RECT 9.455 0.265 9.59 0.33 ;
      RECT 9.08 0.265 9.145 1.14 ;
      RECT 9.32 0.49 9.385 0.625 ;
      RECT 9.08 0.525 9.385 0.59 ;
      RECT 8.935 0.265 9 1.14 ;
      RECT 8.865 0.9775 9 1.0425 ;
      RECT 7.68 0.265 7.745 1.14 ;
      RECT 7.61 0.265 7.745 0.33 ;
      RECT 7.42 0.265 7.485 1.14 ;
      RECT 7.3475 0.265 7.485 0.33 ;
      RECT 7.16 0.265 7.225 1.14 ;
      RECT 7.16 0.625 7.355 0.69 ;
      RECT 7.015 0.265 7.08 1.14 ;
      RECT 6.885 0.9775 7.08 1.0425 ;
      RECT 6.755 0.265 6.82 1.14 ;
      RECT 6.755 0.265 6.89 0.33 ;
      RECT 6.38 0.265 6.445 1.14 ;
      RECT 6.62 0.49 6.685 0.625 ;
      RECT 6.38 0.525 6.685 0.59 ;
      RECT 6.235 0.265 6.3 1.14 ;
      RECT 6.165 0.9775 6.3 1.0425 ;
      RECT 4.98 0.265 5.045 1.14 ;
      RECT 4.91 0.265 5.045 0.33 ;
      RECT 4.72 0.265 4.785 1.14 ;
      RECT 4.6475 0.265 4.785 0.33 ;
      RECT 4.46 0.265 4.525 1.14 ;
      RECT 4.46 0.625 4.655 0.69 ;
      RECT 4.315 0.265 4.38 1.14 ;
      RECT 4.185 0.9775 4.38 1.0425 ;
      RECT 4.055 0.265 4.12 1.14 ;
      RECT 4.055 0.265 4.19 0.33 ;
      RECT 3.68 0.265 3.745 1.14 ;
      RECT 3.92 0.49 3.985 0.625 ;
      RECT 3.68 0.525 3.985 0.59 ;
      RECT 3.535 0.265 3.6 1.14 ;
      RECT 3.465 0.9775 3.6 1.0425 ;
      RECT 2.28 0.265 2.345 1.14 ;
      RECT 2.21 0.265 2.345 0.33 ;
      RECT 2.02 0.265 2.085 1.14 ;
      RECT 1.9475 0.265 2.085 0.33 ;
      RECT 1.76 0.265 1.825 1.14 ;
      RECT 1.76 0.625 1.955 0.69 ;
      RECT 1.615 0.265 1.68 1.14 ;
      RECT 1.485 0.9775 1.68 1.0425 ;
      RECT 1.355 0.265 1.42 1.14 ;
      RECT 1.355 0.265 1.49 0.33 ;
      RECT 0.98 0.265 1.045 1.14 ;
      RECT 1.22 0.49 1.285 0.625 ;
      RECT 0.98 0.525 1.285 0.59 ;
      RECT 0.835 0.265 0.9 1.14 ;
      RECT 0.765 0.9775 0.9 1.0425 ;
      RECT 88.6575 0.41 88.7225 0.545 ;
      RECT 88.5525 0.77 88.6175 0.905 ;
      RECT 88.4225 0.265 88.4875 1.14 ;
      RECT 87.7725 0.41 87.8375 0.545 ;
      RECT 87.7725 0.77 87.8375 0.905 ;
      RECT 87.6425 0.265 87.7075 1.14 ;
      RECT 87.4425 0.6275 87.5775 0.6925 ;
      RECT 86.9375 0.265 87.0025 1.14 ;
      RECT 86.66 0.41 86.725 0.545 ;
      RECT 86.555 0.77 86.62 0.905 ;
      RECT 86.425 0.265 86.49 1.14 ;
      RECT 85.775 0.41 85.84 0.545 ;
      RECT 85.775 0.77 85.84 0.905 ;
      RECT 85.645 0.265 85.71 1.14 ;
      RECT 85.445 0.6275 85.58 0.6925 ;
      RECT 84.94 0.265 85.005 1.14 ;
      RECT 84.665 0.77 84.73 0.905 ;
      RECT 84.405 0.77 84.47 0.905 ;
      RECT 84.13 0.265 84.195 1.14 ;
      RECT 83.755 0.265 83.82 1.14 ;
      RECT 83.61 0.265 83.675 1.14 ;
      RECT 83.15 0.77 83.215 0.905 ;
      RECT 82.89 0.77 82.955 0.905 ;
      RECT 82.485 0.565 82.55 0.7 ;
      RECT 82.11 0.69 82.175 0.825 ;
      RECT 81.705 0.77 81.77 0.905 ;
      RECT 81.43 0.265 81.495 1.14 ;
      RECT 81.055 0.265 81.12 1.14 ;
      RECT 80.91 0.265 80.975 1.14 ;
      RECT 80.45 0.77 80.515 0.905 ;
      RECT 80.19 0.77 80.255 0.905 ;
      RECT 79.785 0.565 79.85 0.7 ;
      RECT 79.41 0.69 79.475 0.825 ;
      RECT 79.005 0.77 79.07 0.905 ;
      RECT 78.73 0.265 78.795 1.14 ;
      RECT 78.355 0.265 78.42 1.14 ;
      RECT 78.21 0.265 78.275 1.14 ;
      RECT 77.75 0.77 77.815 0.905 ;
      RECT 77.49 0.77 77.555 0.905 ;
      RECT 77.085 0.565 77.15 0.7 ;
      RECT 76.71 0.69 76.775 0.825 ;
      RECT 76.305 0.77 76.37 0.905 ;
      RECT 76.03 0.265 76.095 1.14 ;
      RECT 75.655 0.265 75.72 1.14 ;
      RECT 75.51 0.265 75.575 1.14 ;
      RECT 75.05 0.77 75.115 0.905 ;
      RECT 74.79 0.77 74.855 0.905 ;
      RECT 74.385 0.565 74.45 0.7 ;
      RECT 74.01 0.69 74.075 0.825 ;
      RECT 73.605 0.77 73.67 0.905 ;
      RECT 73.33 0.265 73.395 1.14 ;
      RECT 72.955 0.265 73.02 1.14 ;
      RECT 72.81 0.265 72.875 1.14 ;
      RECT 72.35 0.77 72.415 0.905 ;
      RECT 72.09 0.77 72.155 0.905 ;
      RECT 71.685 0.565 71.75 0.7 ;
      RECT 71.31 0.69 71.375 0.825 ;
      RECT 70.905 0.77 70.97 0.905 ;
      RECT 70.63 0.265 70.695 1.14 ;
      RECT 70.255 0.265 70.32 1.14 ;
      RECT 70.11 0.265 70.175 1.14 ;
      RECT 69.65 0.77 69.715 0.905 ;
      RECT 69.39 0.77 69.455 0.905 ;
      RECT 68.985 0.565 69.05 0.7 ;
      RECT 68.61 0.69 68.675 0.825 ;
      RECT 68.205 0.77 68.27 0.905 ;
      RECT 67.93 0.265 67.995 1.14 ;
      RECT 67.555 0.265 67.62 1.14 ;
      RECT 67.41 0.265 67.475 1.14 ;
      RECT 66.95 0.77 67.015 0.905 ;
      RECT 66.69 0.77 66.755 0.905 ;
      RECT 66.285 0.565 66.35 0.7 ;
      RECT 65.91 0.69 65.975 0.825 ;
      RECT 65.505 0.77 65.57 0.905 ;
      RECT 65.23 0.265 65.295 1.14 ;
      RECT 64.855 0.265 64.92 1.14 ;
      RECT 64.71 0.265 64.775 1.14 ;
      RECT 64.25 0.77 64.315 0.905 ;
      RECT 63.99 0.77 64.055 0.905 ;
      RECT 63.585 0.565 63.65 0.7 ;
      RECT 63.21 0.69 63.275 0.825 ;
      RECT 62.805 0.77 62.87 0.905 ;
      RECT 62.53 0.265 62.595 1.14 ;
      RECT 62.155 0.265 62.22 1.14 ;
      RECT 62.01 0.265 62.075 1.14 ;
      RECT 61.55 0.77 61.615 0.905 ;
      RECT 61.29 0.77 61.355 0.905 ;
      RECT 60.885 0.565 60.95 0.7 ;
      RECT 60.51 0.69 60.575 0.825 ;
      RECT 60.105 0.77 60.17 0.905 ;
      RECT 59.83 0.265 59.895 1.14 ;
      RECT 59.455 0.265 59.52 1.14 ;
      RECT 59.31 0.265 59.375 1.14 ;
      RECT 58.85 0.77 58.915 0.905 ;
      RECT 58.59 0.77 58.655 0.905 ;
      RECT 58.185 0.565 58.25 0.7 ;
      RECT 57.81 0.69 57.875 0.825 ;
      RECT 57.405 0.77 57.47 0.905 ;
      RECT 57.13 0.265 57.195 1.14 ;
      RECT 56.755 0.265 56.82 1.14 ;
      RECT 56.61 0.265 56.675 1.14 ;
      RECT 56.15 0.77 56.215 0.905 ;
      RECT 55.89 0.77 55.955 0.905 ;
      RECT 55.485 0.565 55.55 0.7 ;
      RECT 55.11 0.69 55.175 0.825 ;
      RECT 54.705 0.77 54.77 0.905 ;
      RECT 54.43 0.265 54.495 1.14 ;
      RECT 54.055 0.265 54.12 1.14 ;
      RECT 53.91 0.265 53.975 1.14 ;
      RECT 53.45 0.77 53.515 0.905 ;
      RECT 53.19 0.77 53.255 0.905 ;
      RECT 52.785 0.565 52.85 0.7 ;
      RECT 52.41 0.69 52.475 0.825 ;
      RECT 52.005 0.77 52.07 0.905 ;
      RECT 51.73 0.265 51.795 1.14 ;
      RECT 51.355 0.265 51.42 1.14 ;
      RECT 51.21 0.265 51.275 1.14 ;
      RECT 50.75 0.77 50.815 0.905 ;
      RECT 50.49 0.77 50.555 0.905 ;
      RECT 50.085 0.565 50.15 0.7 ;
      RECT 49.71 0.69 49.775 0.825 ;
      RECT 49.305 0.77 49.37 0.905 ;
      RECT 49.03 0.265 49.095 1.14 ;
      RECT 48.655 0.265 48.72 1.14 ;
      RECT 48.51 0.265 48.575 1.14 ;
      RECT 48.05 0.77 48.115 0.905 ;
      RECT 47.79 0.77 47.855 0.905 ;
      RECT 47.385 0.565 47.45 0.7 ;
      RECT 47.01 0.69 47.075 0.825 ;
      RECT 46.605 0.77 46.67 0.905 ;
      RECT 46.33 0.265 46.395 1.14 ;
      RECT 45.955 0.265 46.02 1.14 ;
      RECT 45.81 0.265 45.875 1.14 ;
      RECT 45.35 0.77 45.415 0.905 ;
      RECT 45.09 0.77 45.155 0.905 ;
      RECT 44.685 0.565 44.75 0.7 ;
      RECT 44.31 0.69 44.375 0.825 ;
      RECT 43.905 0.77 43.97 0.905 ;
      RECT 43.63 0.265 43.695 1.14 ;
      RECT 43.255 0.265 43.32 1.14 ;
      RECT 43.11 0.265 43.175 1.14 ;
      RECT 42.65 0.77 42.715 0.905 ;
      RECT 42.39 0.77 42.455 0.905 ;
      RECT 41.985 0.565 42.05 0.7 ;
      RECT 41.61 0.69 41.675 0.825 ;
      RECT 41.205 0.77 41.27 0.905 ;
      RECT 40.93 0.265 40.995 1.14 ;
      RECT 40.555 0.265 40.62 1.14 ;
      RECT 40.41 0.265 40.475 1.14 ;
      RECT 39.95 0.77 40.015 0.905 ;
      RECT 39.69 0.77 39.755 0.905 ;
      RECT 39.285 0.565 39.35 0.7 ;
      RECT 38.91 0.69 38.975 0.825 ;
      RECT 38.505 0.77 38.57 0.905 ;
      RECT 38.23 0.265 38.295 1.14 ;
      RECT 37.855 0.265 37.92 1.14 ;
      RECT 37.71 0.265 37.775 1.14 ;
      RECT 37.25 0.77 37.315 0.905 ;
      RECT 36.99 0.77 37.055 0.905 ;
      RECT 36.585 0.565 36.65 0.7 ;
      RECT 36.21 0.69 36.275 0.825 ;
      RECT 35.805 0.77 35.87 0.905 ;
      RECT 35.53 0.265 35.595 1.14 ;
      RECT 35.155 0.265 35.22 1.14 ;
      RECT 35.01 0.265 35.075 1.14 ;
      RECT 34.55 0.77 34.615 0.905 ;
      RECT 34.29 0.77 34.355 0.905 ;
      RECT 33.885 0.565 33.95 0.7 ;
      RECT 33.51 0.69 33.575 0.825 ;
      RECT 33.105 0.77 33.17 0.905 ;
      RECT 32.83 0.265 32.895 1.14 ;
      RECT 32.455 0.265 32.52 1.14 ;
      RECT 32.31 0.265 32.375 1.14 ;
      RECT 31.85 0.77 31.915 0.905 ;
      RECT 31.59 0.77 31.655 0.905 ;
      RECT 31.185 0.565 31.25 0.7 ;
      RECT 30.81 0.69 30.875 0.825 ;
      RECT 30.405 0.77 30.47 0.905 ;
      RECT 30.13 0.265 30.195 1.14 ;
      RECT 29.755 0.265 29.82 1.14 ;
      RECT 29.61 0.265 29.675 1.14 ;
      RECT 29.15 0.77 29.215 0.905 ;
      RECT 28.89 0.77 28.955 0.905 ;
      RECT 28.485 0.565 28.55 0.7 ;
      RECT 28.11 0.69 28.175 0.825 ;
      RECT 27.705 0.77 27.77 0.905 ;
      RECT 27.43 0.265 27.495 1.14 ;
      RECT 27.055 0.265 27.12 1.14 ;
      RECT 26.91 0.265 26.975 1.14 ;
      RECT 26.45 0.77 26.515 0.905 ;
      RECT 26.19 0.77 26.255 0.905 ;
      RECT 25.785 0.565 25.85 0.7 ;
      RECT 25.41 0.69 25.475 0.825 ;
      RECT 25.005 0.77 25.07 0.905 ;
      RECT 24.73 0.265 24.795 1.14 ;
      RECT 24.355 0.265 24.42 1.14 ;
      RECT 24.21 0.265 24.275 1.14 ;
      RECT 23.75 0.77 23.815 0.905 ;
      RECT 23.49 0.77 23.555 0.905 ;
      RECT 23.085 0.565 23.15 0.7 ;
      RECT 22.71 0.69 22.775 0.825 ;
      RECT 22.305 0.77 22.37 0.905 ;
      RECT 22.03 0.265 22.095 1.14 ;
      RECT 21.655 0.265 21.72 1.14 ;
      RECT 21.51 0.265 21.575 1.14 ;
      RECT 21.05 0.77 21.115 0.905 ;
      RECT 20.79 0.77 20.855 0.905 ;
      RECT 20.385 0.565 20.45 0.7 ;
      RECT 20.01 0.69 20.075 0.825 ;
      RECT 19.605 0.77 19.67 0.905 ;
      RECT 19.33 0.265 19.395 1.14 ;
      RECT 18.955 0.265 19.02 1.14 ;
      RECT 18.81 0.265 18.875 1.14 ;
      RECT 18.35 0.77 18.415 0.905 ;
      RECT 18.09 0.77 18.155 0.905 ;
      RECT 17.685 0.565 17.75 0.7 ;
      RECT 17.31 0.69 17.375 0.825 ;
      RECT 16.905 0.77 16.97 0.905 ;
      RECT 16.63 0.265 16.695 1.14 ;
      RECT 16.255 0.265 16.32 1.14 ;
      RECT 16.11 0.265 16.175 1.14 ;
      RECT 15.65 0.77 15.715 0.905 ;
      RECT 15.39 0.77 15.455 0.905 ;
      RECT 14.985 0.565 15.05 0.7 ;
      RECT 14.61 0.69 14.675 0.825 ;
      RECT 14.205 0.77 14.27 0.905 ;
      RECT 13.93 0.265 13.995 1.14 ;
      RECT 13.555 0.265 13.62 1.14 ;
      RECT 13.41 0.265 13.475 1.14 ;
      RECT 12.95 0.77 13.015 0.905 ;
      RECT 12.69 0.77 12.755 0.905 ;
      RECT 12.285 0.565 12.35 0.7 ;
      RECT 11.91 0.69 11.975 0.825 ;
      RECT 11.505 0.77 11.57 0.905 ;
      RECT 11.23 0.265 11.295 1.14 ;
      RECT 10.855 0.265 10.92 1.14 ;
      RECT 10.71 0.265 10.775 1.14 ;
      RECT 10.25 0.77 10.315 0.905 ;
      RECT 9.99 0.77 10.055 0.905 ;
      RECT 9.585 0.565 9.65 0.7 ;
      RECT 9.21 0.69 9.275 0.825 ;
      RECT 8.805 0.77 8.87 0.905 ;
      RECT 8.53 0.265 8.595 1.14 ;
      RECT 8.155 0.265 8.22 1.14 ;
      RECT 8.01 0.265 8.075 1.14 ;
      RECT 7.55 0.77 7.615 0.905 ;
      RECT 7.29 0.77 7.355 0.905 ;
      RECT 6.885 0.565 6.95 0.7 ;
      RECT 6.51 0.69 6.575 0.825 ;
      RECT 6.105 0.77 6.17 0.905 ;
      RECT 5.83 0.265 5.895 1.14 ;
      RECT 5.455 0.265 5.52 1.14 ;
      RECT 5.31 0.265 5.375 1.14 ;
      RECT 4.85 0.77 4.915 0.905 ;
      RECT 4.59 0.77 4.655 0.905 ;
      RECT 4.185 0.565 4.25 0.7 ;
      RECT 3.81 0.69 3.875 0.825 ;
      RECT 3.405 0.77 3.47 0.905 ;
      RECT 3.13 0.265 3.195 1.14 ;
      RECT 2.755 0.265 2.82 1.14 ;
      RECT 2.61 0.265 2.675 1.14 ;
      RECT 2.15 0.77 2.215 0.905 ;
      RECT 1.89 0.77 1.955 0.905 ;
      RECT 1.485 0.565 1.55 0.7 ;
      RECT 1.11 0.69 1.175 0.825 ;
      RECT 0.705 0.77 0.77 0.905 ;
      RECT 0.43 0.265 0.495 1.14 ;
      RECT 0.055 0.265 0.12 1.14 ;
    LAYER metal2 ;
      RECT 88.795 0.5825 88.865 0.7175 ;
      RECT 87.91 0.5825 87.98 0.7175 ;
      RECT 87.91 0.615 88.865 0.685 ;
      RECT 88.1925 0.5575 88.3275 0.685 ;
      RECT 88.655 0.41 88.725 0.545 ;
      RECT 87.77 0.41 87.84 0.545 ;
      RECT 86.935 0.41 87.005 0.545 ;
      RECT 86.935 0.41 88.725 0.48 ;
      RECT 88.55 0.77 88.62 0.905 ;
      RECT 87.77 0.77 87.84 0.905 ;
      RECT 87.31 0.77 87.38 0.905 ;
      RECT 87.31 0.8025 88.62 0.8725 ;
      RECT 87.4425 0.6225 87.5775 0.695 ;
      RECT 87.4425 0.6225 87.5825 0.6925 ;
      RECT 86.7975 0.5825 86.8675 0.7175 ;
      RECT 85.9125 0.5825 85.9825 0.7175 ;
      RECT 85.9125 0.615 86.8675 0.685 ;
      RECT 86.195 0.5575 86.33 0.685 ;
      RECT 86.6575 0.41 86.7275 0.545 ;
      RECT 85.7725 0.41 85.8425 0.545 ;
      RECT 84.9375 0.41 85.0075 0.545 ;
      RECT 84.9375 0.41 86.7275 0.48 ;
      RECT 86.5525 0.77 86.6225 0.905 ;
      RECT 85.7725 0.77 85.8425 0.905 ;
      RECT 85.3125 0.77 85.3825 0.905 ;
      RECT 85.3125 0.8025 86.6225 0.8725 ;
      RECT 85.445 0.6225 85.58 0.695 ;
      RECT 85.445 0.6225 85.585 0.6925 ;
      RECT 84.725 0.255 84.86 0.3325 ;
      RECT 84.7225 0.255 84.8625 0.325 ;
      RECT 83.7525 0.9475 83.8225 1.0825 ;
      RECT 83.7525 0.98 84.7325 1.05 ;
      RECT 84.6625 0.77 84.7325 1.05 ;
      RECT 84.4025 0.77 84.4725 0.905 ;
      RECT 84.1275 0.77 84.1975 0.905 ;
      RECT 84.1275 0.8025 84.4725 0.8725 ;
      RECT 83.6075 0.77 83.6775 0.905 ;
      RECT 83.1475 0.77 83.2175 0.905 ;
      RECT 83.1475 0.8025 83.6775 0.8725 ;
      RECT 83.21 0.255 83.345 0.3325 ;
      RECT 83.2075 0.255 83.3475 0.325 ;
      RECT 81.4275 1.255 82.9575 1.325 ;
      RECT 82.8875 0.77 82.9575 1.325 ;
      RECT 81.4275 1.005 81.4975 1.325 ;
      RECT 81.5775 1.115 82.76 1.185 ;
      RECT 82.69 0.835 82.76 1.185 ;
      RECT 81.5775 0.835 81.6475 1.185 ;
      RECT 81.0525 0.835 81.1225 1.03 ;
      RECT 82.6225 0.63 82.6925 0.905 ;
      RECT 81.0525 0.835 81.7725 0.905 ;
      RECT 81.7025 0.77 81.7725 0.905 ;
      RECT 82.4825 0.63 82.6925 0.7 ;
      RECT 82.4825 0.565 82.5525 0.7 ;
      RECT 81.765 0.975 82.62 1.045 ;
      RECT 82.1075 0.69 82.1775 1.045 ;
      RECT 80.9075 0.77 80.9775 0.905 ;
      RECT 80.4475 0.77 80.5175 0.905 ;
      RECT 80.4475 0.8025 80.9775 0.8725 ;
      RECT 80.51 0.255 80.645 0.3325 ;
      RECT 80.5075 0.255 80.6475 0.325 ;
      RECT 78.7275 1.255 80.2575 1.325 ;
      RECT 80.1875 0.77 80.2575 1.325 ;
      RECT 78.7275 1.005 78.7975 1.325 ;
      RECT 78.8775 1.115 80.06 1.185 ;
      RECT 79.99 0.835 80.06 1.185 ;
      RECT 78.8775 0.835 78.9475 1.185 ;
      RECT 78.3525 0.835 78.4225 1.03 ;
      RECT 79.9225 0.63 79.9925 0.905 ;
      RECT 78.3525 0.835 79.0725 0.905 ;
      RECT 79.0025 0.77 79.0725 0.905 ;
      RECT 79.7825 0.63 79.9925 0.7 ;
      RECT 79.7825 0.565 79.8525 0.7 ;
      RECT 79.065 0.975 79.92 1.045 ;
      RECT 79.4075 0.69 79.4775 1.045 ;
      RECT 78.2075 0.77 78.2775 0.905 ;
      RECT 77.7475 0.77 77.8175 0.905 ;
      RECT 77.7475 0.8025 78.2775 0.8725 ;
      RECT 77.81 0.255 77.945 0.3325 ;
      RECT 77.8075 0.255 77.9475 0.325 ;
      RECT 76.0275 1.255 77.5575 1.325 ;
      RECT 77.4875 0.77 77.5575 1.325 ;
      RECT 76.0275 1.005 76.0975 1.325 ;
      RECT 76.1775 1.115 77.36 1.185 ;
      RECT 77.29 0.835 77.36 1.185 ;
      RECT 76.1775 0.835 76.2475 1.185 ;
      RECT 75.6525 0.835 75.7225 1.03 ;
      RECT 77.2225 0.63 77.2925 0.905 ;
      RECT 75.6525 0.835 76.3725 0.905 ;
      RECT 76.3025 0.77 76.3725 0.905 ;
      RECT 77.0825 0.63 77.2925 0.7 ;
      RECT 77.0825 0.565 77.1525 0.7 ;
      RECT 76.365 0.975 77.22 1.045 ;
      RECT 76.7075 0.69 76.7775 1.045 ;
      RECT 75.5075 0.77 75.5775 0.905 ;
      RECT 75.0475 0.77 75.1175 0.905 ;
      RECT 75.0475 0.8025 75.5775 0.8725 ;
      RECT 75.11 0.255 75.245 0.3325 ;
      RECT 75.1075 0.255 75.2475 0.325 ;
      RECT 73.3275 1.255 74.8575 1.325 ;
      RECT 74.7875 0.77 74.8575 1.325 ;
      RECT 73.3275 1.005 73.3975 1.325 ;
      RECT 73.4775 1.115 74.66 1.185 ;
      RECT 74.59 0.835 74.66 1.185 ;
      RECT 73.4775 0.835 73.5475 1.185 ;
      RECT 72.9525 0.835 73.0225 1.03 ;
      RECT 74.5225 0.63 74.5925 0.905 ;
      RECT 72.9525 0.835 73.6725 0.905 ;
      RECT 73.6025 0.77 73.6725 0.905 ;
      RECT 74.3825 0.63 74.5925 0.7 ;
      RECT 74.3825 0.565 74.4525 0.7 ;
      RECT 73.665 0.975 74.52 1.045 ;
      RECT 74.0075 0.69 74.0775 1.045 ;
      RECT 72.8075 0.77 72.8775 0.905 ;
      RECT 72.3475 0.77 72.4175 0.905 ;
      RECT 72.3475 0.8025 72.8775 0.8725 ;
      RECT 72.41 0.255 72.545 0.3325 ;
      RECT 72.4075 0.255 72.5475 0.325 ;
      RECT 70.6275 1.255 72.1575 1.325 ;
      RECT 72.0875 0.77 72.1575 1.325 ;
      RECT 70.6275 1.005 70.6975 1.325 ;
      RECT 70.7775 1.115 71.96 1.185 ;
      RECT 71.89 0.835 71.96 1.185 ;
      RECT 70.7775 0.835 70.8475 1.185 ;
      RECT 70.2525 0.835 70.3225 1.03 ;
      RECT 71.8225 0.63 71.8925 0.905 ;
      RECT 70.2525 0.835 70.9725 0.905 ;
      RECT 70.9025 0.77 70.9725 0.905 ;
      RECT 71.6825 0.63 71.8925 0.7 ;
      RECT 71.6825 0.565 71.7525 0.7 ;
      RECT 70.965 0.975 71.82 1.045 ;
      RECT 71.3075 0.69 71.3775 1.045 ;
      RECT 70.1075 0.77 70.1775 0.905 ;
      RECT 69.6475 0.77 69.7175 0.905 ;
      RECT 69.6475 0.8025 70.1775 0.8725 ;
      RECT 69.71 0.255 69.845 0.3325 ;
      RECT 69.7075 0.255 69.8475 0.325 ;
      RECT 67.9275 1.255 69.4575 1.325 ;
      RECT 69.3875 0.77 69.4575 1.325 ;
      RECT 67.9275 1.005 67.9975 1.325 ;
      RECT 68.0775 1.115 69.26 1.185 ;
      RECT 69.19 0.835 69.26 1.185 ;
      RECT 68.0775 0.835 68.1475 1.185 ;
      RECT 67.5525 0.835 67.6225 1.03 ;
      RECT 69.1225 0.63 69.1925 0.905 ;
      RECT 67.5525 0.835 68.2725 0.905 ;
      RECT 68.2025 0.77 68.2725 0.905 ;
      RECT 68.9825 0.63 69.1925 0.7 ;
      RECT 68.9825 0.565 69.0525 0.7 ;
      RECT 68.265 0.975 69.12 1.045 ;
      RECT 68.6075 0.69 68.6775 1.045 ;
      RECT 67.4075 0.77 67.4775 0.905 ;
      RECT 66.9475 0.77 67.0175 0.905 ;
      RECT 66.9475 0.8025 67.4775 0.8725 ;
      RECT 67.01 0.255 67.145 0.3325 ;
      RECT 67.0075 0.255 67.1475 0.325 ;
      RECT 65.2275 1.255 66.7575 1.325 ;
      RECT 66.6875 0.77 66.7575 1.325 ;
      RECT 65.2275 1.005 65.2975 1.325 ;
      RECT 65.3775 1.115 66.56 1.185 ;
      RECT 66.49 0.835 66.56 1.185 ;
      RECT 65.3775 0.835 65.4475 1.185 ;
      RECT 64.8525 0.835 64.9225 1.03 ;
      RECT 66.4225 0.63 66.4925 0.905 ;
      RECT 64.8525 0.835 65.5725 0.905 ;
      RECT 65.5025 0.77 65.5725 0.905 ;
      RECT 66.2825 0.63 66.4925 0.7 ;
      RECT 66.2825 0.565 66.3525 0.7 ;
      RECT 65.565 0.975 66.42 1.045 ;
      RECT 65.9075 0.69 65.9775 1.045 ;
      RECT 64.7075 0.77 64.7775 0.905 ;
      RECT 64.2475 0.77 64.3175 0.905 ;
      RECT 64.2475 0.8025 64.7775 0.8725 ;
      RECT 64.31 0.255 64.445 0.3325 ;
      RECT 64.3075 0.255 64.4475 0.325 ;
      RECT 62.5275 1.255 64.0575 1.325 ;
      RECT 63.9875 0.77 64.0575 1.325 ;
      RECT 62.5275 1.005 62.5975 1.325 ;
      RECT 62.6775 1.115 63.86 1.185 ;
      RECT 63.79 0.835 63.86 1.185 ;
      RECT 62.6775 0.835 62.7475 1.185 ;
      RECT 62.1525 0.835 62.2225 1.03 ;
      RECT 63.7225 0.63 63.7925 0.905 ;
      RECT 62.1525 0.835 62.8725 0.905 ;
      RECT 62.8025 0.77 62.8725 0.905 ;
      RECT 63.5825 0.63 63.7925 0.7 ;
      RECT 63.5825 0.565 63.6525 0.7 ;
      RECT 62.865 0.975 63.72 1.045 ;
      RECT 63.2075 0.69 63.2775 1.045 ;
      RECT 62.0075 0.77 62.0775 0.905 ;
      RECT 61.5475 0.77 61.6175 0.905 ;
      RECT 61.5475 0.8025 62.0775 0.8725 ;
      RECT 61.61 0.255 61.745 0.3325 ;
      RECT 61.6075 0.255 61.7475 0.325 ;
      RECT 59.8275 1.255 61.3575 1.325 ;
      RECT 61.2875 0.77 61.3575 1.325 ;
      RECT 59.8275 1.005 59.8975 1.325 ;
      RECT 59.9775 1.115 61.16 1.185 ;
      RECT 61.09 0.835 61.16 1.185 ;
      RECT 59.9775 0.835 60.0475 1.185 ;
      RECT 59.4525 0.835 59.5225 1.03 ;
      RECT 61.0225 0.63 61.0925 0.905 ;
      RECT 59.4525 0.835 60.1725 0.905 ;
      RECT 60.1025 0.77 60.1725 0.905 ;
      RECT 60.8825 0.63 61.0925 0.7 ;
      RECT 60.8825 0.565 60.9525 0.7 ;
      RECT 60.165 0.975 61.02 1.045 ;
      RECT 60.5075 0.69 60.5775 1.045 ;
      RECT 59.3075 0.77 59.3775 0.905 ;
      RECT 58.8475 0.77 58.9175 0.905 ;
      RECT 58.8475 0.8025 59.3775 0.8725 ;
      RECT 58.91 0.255 59.045 0.3325 ;
      RECT 58.9075 0.255 59.0475 0.325 ;
      RECT 57.1275 1.255 58.6575 1.325 ;
      RECT 58.5875 0.77 58.6575 1.325 ;
      RECT 57.1275 1.005 57.1975 1.325 ;
      RECT 57.2775 1.115 58.46 1.185 ;
      RECT 58.39 0.835 58.46 1.185 ;
      RECT 57.2775 0.835 57.3475 1.185 ;
      RECT 56.7525 0.835 56.8225 1.03 ;
      RECT 58.3225 0.63 58.3925 0.905 ;
      RECT 56.7525 0.835 57.4725 0.905 ;
      RECT 57.4025 0.77 57.4725 0.905 ;
      RECT 58.1825 0.63 58.3925 0.7 ;
      RECT 58.1825 0.565 58.2525 0.7 ;
      RECT 57.465 0.975 58.32 1.045 ;
      RECT 57.8075 0.69 57.8775 1.045 ;
      RECT 56.6075 0.77 56.6775 0.905 ;
      RECT 56.1475 0.77 56.2175 0.905 ;
      RECT 56.1475 0.8025 56.6775 0.8725 ;
      RECT 56.21 0.255 56.345 0.3325 ;
      RECT 56.2075 0.255 56.3475 0.325 ;
      RECT 54.4275 1.255 55.9575 1.325 ;
      RECT 55.8875 0.77 55.9575 1.325 ;
      RECT 54.4275 1.005 54.4975 1.325 ;
      RECT 54.5775 1.115 55.76 1.185 ;
      RECT 55.69 0.835 55.76 1.185 ;
      RECT 54.5775 0.835 54.6475 1.185 ;
      RECT 54.0525 0.835 54.1225 1.03 ;
      RECT 55.6225 0.63 55.6925 0.905 ;
      RECT 54.0525 0.835 54.7725 0.905 ;
      RECT 54.7025 0.77 54.7725 0.905 ;
      RECT 55.4825 0.63 55.6925 0.7 ;
      RECT 55.4825 0.565 55.5525 0.7 ;
      RECT 54.765 0.975 55.62 1.045 ;
      RECT 55.1075 0.69 55.1775 1.045 ;
      RECT 53.9075 0.77 53.9775 0.905 ;
      RECT 53.4475 0.77 53.5175 0.905 ;
      RECT 53.4475 0.8025 53.9775 0.8725 ;
      RECT 53.51 0.255 53.645 0.3325 ;
      RECT 53.5075 0.255 53.6475 0.325 ;
      RECT 51.7275 1.255 53.2575 1.325 ;
      RECT 53.1875 0.77 53.2575 1.325 ;
      RECT 51.7275 1.005 51.7975 1.325 ;
      RECT 51.8775 1.115 53.06 1.185 ;
      RECT 52.99 0.835 53.06 1.185 ;
      RECT 51.8775 0.835 51.9475 1.185 ;
      RECT 51.3525 0.835 51.4225 1.03 ;
      RECT 52.9225 0.63 52.9925 0.905 ;
      RECT 51.3525 0.835 52.0725 0.905 ;
      RECT 52.0025 0.77 52.0725 0.905 ;
      RECT 52.7825 0.63 52.9925 0.7 ;
      RECT 52.7825 0.565 52.8525 0.7 ;
      RECT 52.065 0.975 52.92 1.045 ;
      RECT 52.4075 0.69 52.4775 1.045 ;
      RECT 51.2075 0.77 51.2775 0.905 ;
      RECT 50.7475 0.77 50.8175 0.905 ;
      RECT 50.7475 0.8025 51.2775 0.8725 ;
      RECT 50.81 0.255 50.945 0.3325 ;
      RECT 50.8075 0.255 50.9475 0.325 ;
      RECT 49.0275 1.255 50.5575 1.325 ;
      RECT 50.4875 0.77 50.5575 1.325 ;
      RECT 49.0275 1.005 49.0975 1.325 ;
      RECT 49.1775 1.115 50.36 1.185 ;
      RECT 50.29 0.835 50.36 1.185 ;
      RECT 49.1775 0.835 49.2475 1.185 ;
      RECT 48.6525 0.835 48.7225 1.03 ;
      RECT 50.2225 0.63 50.2925 0.905 ;
      RECT 48.6525 0.835 49.3725 0.905 ;
      RECT 49.3025 0.77 49.3725 0.905 ;
      RECT 50.0825 0.63 50.2925 0.7 ;
      RECT 50.0825 0.565 50.1525 0.7 ;
      RECT 49.365 0.975 50.22 1.045 ;
      RECT 49.7075 0.69 49.7775 1.045 ;
      RECT 48.5075 0.77 48.5775 0.905 ;
      RECT 48.0475 0.77 48.1175 0.905 ;
      RECT 48.0475 0.8025 48.5775 0.8725 ;
      RECT 48.11 0.255 48.245 0.3325 ;
      RECT 48.1075 0.255 48.2475 0.325 ;
      RECT 46.3275 1.255 47.8575 1.325 ;
      RECT 47.7875 0.77 47.8575 1.325 ;
      RECT 46.3275 1.005 46.3975 1.325 ;
      RECT 46.4775 1.115 47.66 1.185 ;
      RECT 47.59 0.835 47.66 1.185 ;
      RECT 46.4775 0.835 46.5475 1.185 ;
      RECT 45.9525 0.835 46.0225 1.03 ;
      RECT 47.5225 0.63 47.5925 0.905 ;
      RECT 45.9525 0.835 46.6725 0.905 ;
      RECT 46.6025 0.77 46.6725 0.905 ;
      RECT 47.3825 0.63 47.5925 0.7 ;
      RECT 47.3825 0.565 47.4525 0.7 ;
      RECT 46.665 0.975 47.52 1.045 ;
      RECT 47.0075 0.69 47.0775 1.045 ;
      RECT 45.8075 0.77 45.8775 0.905 ;
      RECT 45.3475 0.77 45.4175 0.905 ;
      RECT 45.3475 0.8025 45.8775 0.8725 ;
      RECT 45.41 0.255 45.545 0.3325 ;
      RECT 45.4075 0.255 45.5475 0.325 ;
      RECT 43.6275 1.255 45.1575 1.325 ;
      RECT 45.0875 0.77 45.1575 1.325 ;
      RECT 43.6275 1.005 43.6975 1.325 ;
      RECT 43.7775 1.115 44.96 1.185 ;
      RECT 44.89 0.835 44.96 1.185 ;
      RECT 43.7775 0.835 43.8475 1.185 ;
      RECT 43.2525 0.835 43.3225 1.03 ;
      RECT 44.8225 0.63 44.8925 0.905 ;
      RECT 43.2525 0.835 43.9725 0.905 ;
      RECT 43.9025 0.77 43.9725 0.905 ;
      RECT 44.6825 0.63 44.8925 0.7 ;
      RECT 44.6825 0.565 44.7525 0.7 ;
      RECT 43.965 0.975 44.82 1.045 ;
      RECT 44.3075 0.69 44.3775 1.045 ;
      RECT 43.1075 0.77 43.1775 0.905 ;
      RECT 42.6475 0.77 42.7175 0.905 ;
      RECT 42.6475 0.8025 43.1775 0.8725 ;
      RECT 42.71 0.255 42.845 0.3325 ;
      RECT 42.7075 0.255 42.8475 0.325 ;
      RECT 40.9275 1.255 42.4575 1.325 ;
      RECT 42.3875 0.77 42.4575 1.325 ;
      RECT 40.9275 1.005 40.9975 1.325 ;
      RECT 41.0775 1.115 42.26 1.185 ;
      RECT 42.19 0.835 42.26 1.185 ;
      RECT 41.0775 0.835 41.1475 1.185 ;
      RECT 40.5525 0.835 40.6225 1.03 ;
      RECT 42.1225 0.63 42.1925 0.905 ;
      RECT 40.5525 0.835 41.2725 0.905 ;
      RECT 41.2025 0.77 41.2725 0.905 ;
      RECT 41.9825 0.63 42.1925 0.7 ;
      RECT 41.9825 0.565 42.0525 0.7 ;
      RECT 41.265 0.975 42.12 1.045 ;
      RECT 41.6075 0.69 41.6775 1.045 ;
      RECT 40.4075 0.77 40.4775 0.905 ;
      RECT 39.9475 0.77 40.0175 0.905 ;
      RECT 39.9475 0.8025 40.4775 0.8725 ;
      RECT 40.01 0.255 40.145 0.3325 ;
      RECT 40.0075 0.255 40.1475 0.325 ;
      RECT 38.2275 1.255 39.7575 1.325 ;
      RECT 39.6875 0.77 39.7575 1.325 ;
      RECT 38.2275 1.005 38.2975 1.325 ;
      RECT 38.3775 1.115 39.56 1.185 ;
      RECT 39.49 0.835 39.56 1.185 ;
      RECT 38.3775 0.835 38.4475 1.185 ;
      RECT 37.8525 0.835 37.9225 1.03 ;
      RECT 39.4225 0.63 39.4925 0.905 ;
      RECT 37.8525 0.835 38.5725 0.905 ;
      RECT 38.5025 0.77 38.5725 0.905 ;
      RECT 39.2825 0.63 39.4925 0.7 ;
      RECT 39.2825 0.565 39.3525 0.7 ;
      RECT 38.565 0.975 39.42 1.045 ;
      RECT 38.9075 0.69 38.9775 1.045 ;
      RECT 37.7075 0.77 37.7775 0.905 ;
      RECT 37.2475 0.77 37.3175 0.905 ;
      RECT 37.2475 0.8025 37.7775 0.8725 ;
      RECT 37.31 0.255 37.445 0.3325 ;
      RECT 37.3075 0.255 37.4475 0.325 ;
      RECT 35.5275 1.255 37.0575 1.325 ;
      RECT 36.9875 0.77 37.0575 1.325 ;
      RECT 35.5275 1.005 35.5975 1.325 ;
      RECT 35.6775 1.115 36.86 1.185 ;
      RECT 36.79 0.835 36.86 1.185 ;
      RECT 35.6775 0.835 35.7475 1.185 ;
      RECT 35.1525 0.835 35.2225 1.03 ;
      RECT 36.7225 0.63 36.7925 0.905 ;
      RECT 35.1525 0.835 35.8725 0.905 ;
      RECT 35.8025 0.77 35.8725 0.905 ;
      RECT 36.5825 0.63 36.7925 0.7 ;
      RECT 36.5825 0.565 36.6525 0.7 ;
      RECT 35.865 0.975 36.72 1.045 ;
      RECT 36.2075 0.69 36.2775 1.045 ;
      RECT 35.0075 0.77 35.0775 0.905 ;
      RECT 34.5475 0.77 34.6175 0.905 ;
      RECT 34.5475 0.8025 35.0775 0.8725 ;
      RECT 34.61 0.255 34.745 0.3325 ;
      RECT 34.6075 0.255 34.7475 0.325 ;
      RECT 32.8275 1.255 34.3575 1.325 ;
      RECT 34.2875 0.77 34.3575 1.325 ;
      RECT 32.8275 1.005 32.8975 1.325 ;
      RECT 32.9775 1.115 34.16 1.185 ;
      RECT 34.09 0.835 34.16 1.185 ;
      RECT 32.9775 0.835 33.0475 1.185 ;
      RECT 32.4525 0.835 32.5225 1.03 ;
      RECT 34.0225 0.63 34.0925 0.905 ;
      RECT 32.4525 0.835 33.1725 0.905 ;
      RECT 33.1025 0.77 33.1725 0.905 ;
      RECT 33.8825 0.63 34.0925 0.7 ;
      RECT 33.8825 0.565 33.9525 0.7 ;
      RECT 33.165 0.975 34.02 1.045 ;
      RECT 33.5075 0.69 33.5775 1.045 ;
      RECT 32.3075 0.77 32.3775 0.905 ;
      RECT 31.8475 0.77 31.9175 0.905 ;
      RECT 31.8475 0.8025 32.3775 0.8725 ;
      RECT 31.91 0.255 32.045 0.3325 ;
      RECT 31.9075 0.255 32.0475 0.325 ;
      RECT 30.1275 1.255 31.6575 1.325 ;
      RECT 31.5875 0.77 31.6575 1.325 ;
      RECT 30.1275 1.005 30.1975 1.325 ;
      RECT 30.2775 1.115 31.46 1.185 ;
      RECT 31.39 0.835 31.46 1.185 ;
      RECT 30.2775 0.835 30.3475 1.185 ;
      RECT 29.7525 0.835 29.8225 1.03 ;
      RECT 31.3225 0.63 31.3925 0.905 ;
      RECT 29.7525 0.835 30.4725 0.905 ;
      RECT 30.4025 0.77 30.4725 0.905 ;
      RECT 31.1825 0.63 31.3925 0.7 ;
      RECT 31.1825 0.565 31.2525 0.7 ;
      RECT 30.465 0.975 31.32 1.045 ;
      RECT 30.8075 0.69 30.8775 1.045 ;
      RECT 29.6075 0.77 29.6775 0.905 ;
      RECT 29.1475 0.77 29.2175 0.905 ;
      RECT 29.1475 0.8025 29.6775 0.8725 ;
      RECT 29.21 0.255 29.345 0.3325 ;
      RECT 29.2075 0.255 29.3475 0.325 ;
      RECT 27.4275 1.255 28.9575 1.325 ;
      RECT 28.8875 0.77 28.9575 1.325 ;
      RECT 27.4275 1.005 27.4975 1.325 ;
      RECT 27.5775 1.115 28.76 1.185 ;
      RECT 28.69 0.835 28.76 1.185 ;
      RECT 27.5775 0.835 27.6475 1.185 ;
      RECT 27.0525 0.835 27.1225 1.03 ;
      RECT 28.6225 0.63 28.6925 0.905 ;
      RECT 27.0525 0.835 27.7725 0.905 ;
      RECT 27.7025 0.77 27.7725 0.905 ;
      RECT 28.4825 0.63 28.6925 0.7 ;
      RECT 28.4825 0.565 28.5525 0.7 ;
      RECT 27.765 0.975 28.62 1.045 ;
      RECT 28.1075 0.69 28.1775 1.045 ;
      RECT 26.9075 0.77 26.9775 0.905 ;
      RECT 26.4475 0.77 26.5175 0.905 ;
      RECT 26.4475 0.8025 26.9775 0.8725 ;
      RECT 26.51 0.255 26.645 0.3325 ;
      RECT 26.5075 0.255 26.6475 0.325 ;
      RECT 24.7275 1.255 26.2575 1.325 ;
      RECT 26.1875 0.77 26.2575 1.325 ;
      RECT 24.7275 1.005 24.7975 1.325 ;
      RECT 24.8775 1.115 26.06 1.185 ;
      RECT 25.99 0.835 26.06 1.185 ;
      RECT 24.8775 0.835 24.9475 1.185 ;
      RECT 24.3525 0.835 24.4225 1.03 ;
      RECT 25.9225 0.63 25.9925 0.905 ;
      RECT 24.3525 0.835 25.0725 0.905 ;
      RECT 25.0025 0.77 25.0725 0.905 ;
      RECT 25.7825 0.63 25.9925 0.7 ;
      RECT 25.7825 0.565 25.8525 0.7 ;
      RECT 25.065 0.975 25.92 1.045 ;
      RECT 25.4075 0.69 25.4775 1.045 ;
      RECT 24.2075 0.77 24.2775 0.905 ;
      RECT 23.7475 0.77 23.8175 0.905 ;
      RECT 23.7475 0.8025 24.2775 0.8725 ;
      RECT 23.81 0.255 23.945 0.3325 ;
      RECT 23.8075 0.255 23.9475 0.325 ;
      RECT 22.0275 1.255 23.5575 1.325 ;
      RECT 23.4875 0.77 23.5575 1.325 ;
      RECT 22.0275 1.005 22.0975 1.325 ;
      RECT 22.1775 1.115 23.36 1.185 ;
      RECT 23.29 0.835 23.36 1.185 ;
      RECT 22.1775 0.835 22.2475 1.185 ;
      RECT 21.6525 0.835 21.7225 1.03 ;
      RECT 23.2225 0.63 23.2925 0.905 ;
      RECT 21.6525 0.835 22.3725 0.905 ;
      RECT 22.3025 0.77 22.3725 0.905 ;
      RECT 23.0825 0.63 23.2925 0.7 ;
      RECT 23.0825 0.565 23.1525 0.7 ;
      RECT 22.365 0.975 23.22 1.045 ;
      RECT 22.7075 0.69 22.7775 1.045 ;
      RECT 21.5075 0.77 21.5775 0.905 ;
      RECT 21.0475 0.77 21.1175 0.905 ;
      RECT 21.0475 0.8025 21.5775 0.8725 ;
      RECT 21.11 0.255 21.245 0.3325 ;
      RECT 21.1075 0.255 21.2475 0.325 ;
      RECT 19.3275 1.255 20.8575 1.325 ;
      RECT 20.7875 0.77 20.8575 1.325 ;
      RECT 19.3275 1.005 19.3975 1.325 ;
      RECT 19.4775 1.115 20.66 1.185 ;
      RECT 20.59 0.835 20.66 1.185 ;
      RECT 19.4775 0.835 19.5475 1.185 ;
      RECT 18.9525 0.835 19.0225 1.03 ;
      RECT 20.5225 0.63 20.5925 0.905 ;
      RECT 18.9525 0.835 19.6725 0.905 ;
      RECT 19.6025 0.77 19.6725 0.905 ;
      RECT 20.3825 0.63 20.5925 0.7 ;
      RECT 20.3825 0.565 20.4525 0.7 ;
      RECT 19.665 0.975 20.52 1.045 ;
      RECT 20.0075 0.69 20.0775 1.045 ;
      RECT 18.8075 0.77 18.8775 0.905 ;
      RECT 18.3475 0.77 18.4175 0.905 ;
      RECT 18.3475 0.8025 18.8775 0.8725 ;
      RECT 18.41 0.255 18.545 0.3325 ;
      RECT 18.4075 0.255 18.5475 0.325 ;
      RECT 16.6275 1.255 18.1575 1.325 ;
      RECT 18.0875 0.77 18.1575 1.325 ;
      RECT 16.6275 1.005 16.6975 1.325 ;
      RECT 16.7775 1.115 17.96 1.185 ;
      RECT 17.89 0.835 17.96 1.185 ;
      RECT 16.7775 0.835 16.8475 1.185 ;
      RECT 16.2525 0.835 16.3225 1.03 ;
      RECT 17.8225 0.63 17.8925 0.905 ;
      RECT 16.2525 0.835 16.9725 0.905 ;
      RECT 16.9025 0.77 16.9725 0.905 ;
      RECT 17.6825 0.63 17.8925 0.7 ;
      RECT 17.6825 0.565 17.7525 0.7 ;
      RECT 16.965 0.975 17.82 1.045 ;
      RECT 17.3075 0.69 17.3775 1.045 ;
      RECT 16.1075 0.77 16.1775 0.905 ;
      RECT 15.6475 0.77 15.7175 0.905 ;
      RECT 15.6475 0.8025 16.1775 0.8725 ;
      RECT 15.71 0.255 15.845 0.3325 ;
      RECT 15.7075 0.255 15.8475 0.325 ;
      RECT 13.9275 1.255 15.4575 1.325 ;
      RECT 15.3875 0.77 15.4575 1.325 ;
      RECT 13.9275 1.005 13.9975 1.325 ;
      RECT 14.0775 1.115 15.26 1.185 ;
      RECT 15.19 0.835 15.26 1.185 ;
      RECT 14.0775 0.835 14.1475 1.185 ;
      RECT 13.5525 0.835 13.6225 1.03 ;
      RECT 15.1225 0.63 15.1925 0.905 ;
      RECT 13.5525 0.835 14.2725 0.905 ;
      RECT 14.2025 0.77 14.2725 0.905 ;
      RECT 14.9825 0.63 15.1925 0.7 ;
      RECT 14.9825 0.565 15.0525 0.7 ;
      RECT 14.265 0.975 15.12 1.045 ;
      RECT 14.6075 0.69 14.6775 1.045 ;
      RECT 13.4075 0.77 13.4775 0.905 ;
      RECT 12.9475 0.77 13.0175 0.905 ;
      RECT 12.9475 0.8025 13.4775 0.8725 ;
      RECT 13.01 0.255 13.145 0.3325 ;
      RECT 13.0075 0.255 13.1475 0.325 ;
      RECT 11.2275 1.255 12.7575 1.325 ;
      RECT 12.6875 0.77 12.7575 1.325 ;
      RECT 11.2275 1.005 11.2975 1.325 ;
      RECT 11.3775 1.115 12.56 1.185 ;
      RECT 12.49 0.835 12.56 1.185 ;
      RECT 11.3775 0.835 11.4475 1.185 ;
      RECT 10.8525 0.835 10.9225 1.03 ;
      RECT 12.4225 0.63 12.4925 0.905 ;
      RECT 10.8525 0.835 11.5725 0.905 ;
      RECT 11.5025 0.77 11.5725 0.905 ;
      RECT 12.2825 0.63 12.4925 0.7 ;
      RECT 12.2825 0.565 12.3525 0.7 ;
      RECT 11.565 0.975 12.42 1.045 ;
      RECT 11.9075 0.69 11.9775 1.045 ;
      RECT 10.7075 0.77 10.7775 0.905 ;
      RECT 10.2475 0.77 10.3175 0.905 ;
      RECT 10.2475 0.8025 10.7775 0.8725 ;
      RECT 10.31 0.255 10.445 0.3325 ;
      RECT 10.3075 0.255 10.4475 0.325 ;
      RECT 8.5275 1.255 10.0575 1.325 ;
      RECT 9.9875 0.77 10.0575 1.325 ;
      RECT 8.5275 1.005 8.5975 1.325 ;
      RECT 8.6775 1.115 9.86 1.185 ;
      RECT 9.79 0.835 9.86 1.185 ;
      RECT 8.6775 0.835 8.7475 1.185 ;
      RECT 8.1525 0.835 8.2225 1.03 ;
      RECT 9.7225 0.63 9.7925 0.905 ;
      RECT 8.1525 0.835 8.8725 0.905 ;
      RECT 8.8025 0.77 8.8725 0.905 ;
      RECT 9.5825 0.63 9.7925 0.7 ;
      RECT 9.5825 0.565 9.6525 0.7 ;
      RECT 8.865 0.975 9.72 1.045 ;
      RECT 9.2075 0.69 9.2775 1.045 ;
      RECT 8.0075 0.77 8.0775 0.905 ;
      RECT 7.5475 0.77 7.6175 0.905 ;
      RECT 7.5475 0.8025 8.0775 0.8725 ;
      RECT 7.61 0.255 7.745 0.3325 ;
      RECT 7.6075 0.255 7.7475 0.325 ;
      RECT 5.8275 1.255 7.3575 1.325 ;
      RECT 7.2875 0.77 7.3575 1.325 ;
      RECT 5.8275 1.005 5.8975 1.325 ;
      RECT 5.9775 1.115 7.16 1.185 ;
      RECT 7.09 0.835 7.16 1.185 ;
      RECT 5.9775 0.835 6.0475 1.185 ;
      RECT 5.4525 0.835 5.5225 1.03 ;
      RECT 7.0225 0.63 7.0925 0.905 ;
      RECT 5.4525 0.835 6.1725 0.905 ;
      RECT 6.1025 0.77 6.1725 0.905 ;
      RECT 6.8825 0.63 7.0925 0.7 ;
      RECT 6.8825 0.565 6.9525 0.7 ;
      RECT 6.165 0.975 7.02 1.045 ;
      RECT 6.5075 0.69 6.5775 1.045 ;
      RECT 5.3075 0.77 5.3775 0.905 ;
      RECT 4.8475 0.77 4.9175 0.905 ;
      RECT 4.8475 0.8025 5.3775 0.8725 ;
      RECT 4.91 0.255 5.045 0.3325 ;
      RECT 4.9075 0.255 5.0475 0.325 ;
      RECT 3.1275 1.255 4.6575 1.325 ;
      RECT 4.5875 0.77 4.6575 1.325 ;
      RECT 3.1275 1.005 3.1975 1.325 ;
      RECT 3.2775 1.115 4.46 1.185 ;
      RECT 4.39 0.835 4.46 1.185 ;
      RECT 3.2775 0.835 3.3475 1.185 ;
      RECT 2.7525 0.835 2.8225 1.03 ;
      RECT 4.3225 0.63 4.3925 0.905 ;
      RECT 2.7525 0.835 3.4725 0.905 ;
      RECT 3.4025 0.77 3.4725 0.905 ;
      RECT 4.1825 0.63 4.3925 0.7 ;
      RECT 4.1825 0.565 4.2525 0.7 ;
      RECT 3.465 0.975 4.32 1.045 ;
      RECT 3.8075 0.69 3.8775 1.045 ;
      RECT 2.6075 0.77 2.6775 0.905 ;
      RECT 2.1475 0.77 2.2175 0.905 ;
      RECT 2.1475 0.8025 2.6775 0.8725 ;
      RECT 2.21 0.255 2.345 0.3325 ;
      RECT 2.2075 0.255 2.3475 0.325 ;
      RECT 0.4275 1.255 1.9575 1.325 ;
      RECT 1.8875 0.77 1.9575 1.325 ;
      RECT 0.4275 1.005 0.4975 1.325 ;
      RECT 0.5775 1.115 1.76 1.185 ;
      RECT 1.69 0.835 1.76 1.185 ;
      RECT 0.5775 0.835 0.6475 1.185 ;
      RECT 0.0525 0.835 0.1225 1.03 ;
      RECT 1.6225 0.63 1.6925 0.905 ;
      RECT 0.0525 0.835 0.7725 0.905 ;
      RECT 0.7025 0.77 0.7725 0.905 ;
      RECT 1.4825 0.63 1.6925 0.7 ;
      RECT 1.4825 0.565 1.5525 0.7 ;
      RECT 0.765 0.975 1.62 1.045 ;
      RECT 1.1075 0.69 1.1775 1.045 ;
      RECT 84.33 0.6225 84.47 0.6925 ;
      RECT 82.355 0.2625 83.0825 0.3325 ;
      RECT 82.8175 0.6225 82.9575 0.6925 ;
      RECT 79.655 0.2625 80.3825 0.3325 ;
      RECT 80.1175 0.6225 80.2575 0.6925 ;
      RECT 76.955 0.2625 77.6825 0.3325 ;
      RECT 77.4175 0.6225 77.5575 0.6925 ;
      RECT 74.255 0.2625 74.9825 0.3325 ;
      RECT 74.7175 0.6225 74.8575 0.6925 ;
      RECT 71.555 0.2625 72.2825 0.3325 ;
      RECT 72.0175 0.6225 72.1575 0.6925 ;
      RECT 68.855 0.2625 69.5825 0.3325 ;
      RECT 69.3175 0.6225 69.4575 0.6925 ;
      RECT 66.155 0.2625 66.8825 0.3325 ;
      RECT 66.6175 0.6225 66.7575 0.6925 ;
      RECT 63.455 0.2625 64.1825 0.3325 ;
      RECT 63.9175 0.6225 64.0575 0.6925 ;
      RECT 60.755 0.2625 61.4825 0.3325 ;
      RECT 61.2175 0.6225 61.3575 0.6925 ;
      RECT 58.055 0.2625 58.7825 0.3325 ;
      RECT 58.5175 0.6225 58.6575 0.6925 ;
      RECT 55.355 0.2625 56.0825 0.3325 ;
      RECT 55.8175 0.6225 55.9575 0.6925 ;
      RECT 52.655 0.2625 53.3825 0.3325 ;
      RECT 53.1175 0.6225 53.2575 0.6925 ;
      RECT 49.955 0.2625 50.6825 0.3325 ;
      RECT 50.4175 0.6225 50.5575 0.6925 ;
      RECT 47.255 0.2625 47.9825 0.3325 ;
      RECT 47.7175 0.6225 47.8575 0.6925 ;
      RECT 44.555 0.2625 45.2825 0.3325 ;
      RECT 45.0175 0.6225 45.1575 0.6925 ;
      RECT 41.855 0.2625 42.5825 0.3325 ;
      RECT 42.3175 0.6225 42.4575 0.6925 ;
      RECT 39.155 0.2625 39.8825 0.3325 ;
      RECT 39.6175 0.6225 39.7575 0.6925 ;
      RECT 36.455 0.2625 37.1825 0.3325 ;
      RECT 36.9175 0.6225 37.0575 0.6925 ;
      RECT 33.755 0.2625 34.4825 0.3325 ;
      RECT 34.2175 0.6225 34.3575 0.6925 ;
      RECT 31.055 0.2625 31.7825 0.3325 ;
      RECT 31.5175 0.6225 31.6575 0.6925 ;
      RECT 28.355 0.2625 29.0825 0.3325 ;
      RECT 28.8175 0.6225 28.9575 0.6925 ;
      RECT 25.655 0.2625 26.3825 0.3325 ;
      RECT 26.1175 0.6225 26.2575 0.6925 ;
      RECT 22.955 0.2625 23.6825 0.3325 ;
      RECT 23.4175 0.6225 23.5575 0.6925 ;
      RECT 20.255 0.2625 20.9825 0.3325 ;
      RECT 20.7175 0.6225 20.8575 0.6925 ;
      RECT 17.555 0.2625 18.2825 0.3325 ;
      RECT 18.0175 0.6225 18.1575 0.6925 ;
      RECT 14.855 0.2625 15.5825 0.3325 ;
      RECT 15.3175 0.6225 15.4575 0.6925 ;
      RECT 12.155 0.2625 12.8825 0.3325 ;
      RECT 12.6175 0.6225 12.7575 0.6925 ;
      RECT 9.455 0.2625 10.1825 0.3325 ;
      RECT 9.9175 0.6225 10.0575 0.6925 ;
      RECT 6.755 0.2625 7.4825 0.3325 ;
      RECT 7.2175 0.6225 7.3575 0.6925 ;
      RECT 4.055 0.2625 4.7825 0.3325 ;
      RECT 4.5175 0.6225 4.6575 0.6925 ;
      RECT 1.355 0.2625 2.0825 0.3325 ;
      RECT 1.8175 0.6225 1.9575 0.6925 ;
    LAYER metal3 ;
      RECT 87.4425 0.6225 87.5825 0.6925 ;
      RECT 87.4425 0.255 87.5125 0.6925 ;
      RECT 2.2075 0.255 87.5125 0.325 ;
      RECT 85.445 0.6225 85.585 0.6925 ;
      RECT 84.33 0.6225 84.47 0.6925 ;
      RECT 82.8175 0.6225 82.9575 0.6925 ;
      RECT 80.1175 0.6225 80.2575 0.6925 ;
      RECT 77.4175 0.6225 77.5575 0.6925 ;
      RECT 74.7175 0.6225 74.8575 0.6925 ;
      RECT 72.0175 0.6225 72.1575 0.6925 ;
      RECT 69.3175 0.6225 69.4575 0.6925 ;
      RECT 66.6175 0.6225 66.7575 0.6925 ;
      RECT 63.9175 0.6225 64.0575 0.6925 ;
      RECT 61.2175 0.6225 61.3575 0.6925 ;
      RECT 58.5175 0.6225 58.6575 0.6925 ;
      RECT 55.8175 0.6225 55.9575 0.6925 ;
      RECT 53.1175 0.6225 53.2575 0.6925 ;
      RECT 50.4175 0.6225 50.5575 0.6925 ;
      RECT 47.7175 0.6225 47.8575 0.6925 ;
      RECT 45.0175 0.6225 45.1575 0.6925 ;
      RECT 42.3175 0.6225 42.4575 0.6925 ;
      RECT 39.6175 0.6225 39.7575 0.6925 ;
      RECT 36.9175 0.6225 37.0575 0.6925 ;
      RECT 34.2175 0.6225 34.3575 0.6925 ;
      RECT 31.5175 0.6225 31.6575 0.6925 ;
      RECT 28.8175 0.6225 28.9575 0.6925 ;
      RECT 26.1175 0.6225 26.2575 0.6925 ;
      RECT 23.4175 0.6225 23.5575 0.6925 ;
      RECT 20.7175 0.6225 20.8575 0.6925 ;
      RECT 18.0175 0.6225 18.1575 0.6925 ;
      RECT 15.3175 0.6225 15.4575 0.6925 ;
      RECT 12.6175 0.6225 12.7575 0.6925 ;
      RECT 9.9175 0.6225 10.0575 0.6925 ;
      RECT 7.2175 0.6225 7.3575 0.6925 ;
      RECT 4.5175 0.6225 4.6575 0.6925 ;
      RECT 1.8175 0.6225 1.9575 0.6925 ;
      RECT 85.445 0.395 85.515 0.6925 ;
      RECT 84.33 0.395 84.4 0.6925 ;
      RECT 82.8175 0.395 82.8875 0.6925 ;
      RECT 80.1175 0.395 80.1875 0.6925 ;
      RECT 77.4175 0.395 77.4875 0.6925 ;
      RECT 74.7175 0.395 74.7875 0.6925 ;
      RECT 72.0175 0.395 72.0875 0.6925 ;
      RECT 69.3175 0.395 69.3875 0.6925 ;
      RECT 66.6175 0.395 66.6875 0.6925 ;
      RECT 63.9175 0.395 63.9875 0.6925 ;
      RECT 61.2175 0.395 61.2875 0.6925 ;
      RECT 58.5175 0.395 58.5875 0.6925 ;
      RECT 55.8175 0.395 55.8875 0.6925 ;
      RECT 53.1175 0.395 53.1875 0.6925 ;
      RECT 50.4175 0.395 50.4875 0.6925 ;
      RECT 47.7175 0.395 47.7875 0.6925 ;
      RECT 45.0175 0.395 45.0875 0.6925 ;
      RECT 42.3175 0.395 42.3875 0.6925 ;
      RECT 39.6175 0.395 39.6875 0.6925 ;
      RECT 36.9175 0.395 36.9875 0.6925 ;
      RECT 34.2175 0.395 34.2875 0.6925 ;
      RECT 31.5175 0.395 31.5875 0.6925 ;
      RECT 28.8175 0.395 28.8875 0.6925 ;
      RECT 26.1175 0.395 26.1875 0.6925 ;
      RECT 23.4175 0.395 23.4875 0.6925 ;
      RECT 20.7175 0.395 20.7875 0.6925 ;
      RECT 18.0175 0.395 18.0875 0.6925 ;
      RECT 15.3175 0.395 15.3875 0.6925 ;
      RECT 12.6175 0.395 12.6875 0.6925 ;
      RECT 9.9175 0.395 9.9875 0.6925 ;
      RECT 7.2175 0.395 7.2875 0.6925 ;
      RECT 4.5175 0.395 4.5875 0.6925 ;
      RECT 1.8175 0.395 1.8875 0.6925 ;
      RECT 1.8175 0.395 85.515 0.465 ;
    LAYER via1 ;
      RECT 88.7975 0.6175 88.8625 0.6825 ;
      RECT 88.6575 0.445 88.7225 0.51 ;
      RECT 88.5525 0.805 88.6175 0.87 ;
      RECT 88.2275 0.56 88.2925 0.625 ;
      RECT 87.9125 0.6175 87.9775 0.6825 ;
      RECT 87.7725 0.445 87.8375 0.51 ;
      RECT 87.7725 0.805 87.8375 0.87 ;
      RECT 87.4775 0.6275 87.5425 0.6925 ;
      RECT 87.3125 0.805 87.3775 0.87 ;
      RECT 86.9375 0.445 87.0025 0.51 ;
      RECT 86.8 0.6175 86.865 0.6825 ;
      RECT 86.66 0.445 86.725 0.51 ;
      RECT 86.555 0.805 86.62 0.87 ;
      RECT 86.23 0.56 86.295 0.625 ;
      RECT 85.915 0.6175 85.98 0.6825 ;
      RECT 85.775 0.445 85.84 0.51 ;
      RECT 85.775 0.805 85.84 0.87 ;
      RECT 85.48 0.6275 85.545 0.6925 ;
      RECT 85.315 0.805 85.38 0.87 ;
      RECT 84.94 0.445 85.005 0.51 ;
      RECT 84.76 0.265 84.825 0.33 ;
      RECT 84.665 0.805 84.73 0.87 ;
      RECT 84.405 0.805 84.47 0.87 ;
      RECT 84.3675 0.625 84.4325 0.69 ;
      RECT 84.13 0.805 84.195 0.87 ;
      RECT 83.755 0.9825 83.82 1.0475 ;
      RECT 83.61 0.805 83.675 0.87 ;
      RECT 83.245 0.265 83.31 0.33 ;
      RECT 83.15 0.805 83.215 0.87 ;
      RECT 82.9825 0.265 83.0475 0.33 ;
      RECT 82.89 0.805 82.955 0.87 ;
      RECT 82.855 0.625 82.92 0.69 ;
      RECT 82.52 0.9775 82.585 1.0425 ;
      RECT 82.485 0.6 82.55 0.665 ;
      RECT 82.39 0.265 82.455 0.33 ;
      RECT 82.11 0.725 82.175 0.79 ;
      RECT 81.8 0.9775 81.865 1.0425 ;
      RECT 81.705 0.805 81.77 0.87 ;
      RECT 81.43 1.04 81.495 1.105 ;
      RECT 81.055 0.93 81.12 0.995 ;
      RECT 80.91 0.805 80.975 0.87 ;
      RECT 80.545 0.265 80.61 0.33 ;
      RECT 80.45 0.805 80.515 0.87 ;
      RECT 80.2825 0.265 80.3475 0.33 ;
      RECT 80.19 0.805 80.255 0.87 ;
      RECT 80.155 0.625 80.22 0.69 ;
      RECT 79.82 0.9775 79.885 1.0425 ;
      RECT 79.785 0.6 79.85 0.665 ;
      RECT 79.69 0.265 79.755 0.33 ;
      RECT 79.41 0.725 79.475 0.79 ;
      RECT 79.1 0.9775 79.165 1.0425 ;
      RECT 79.005 0.805 79.07 0.87 ;
      RECT 78.73 1.04 78.795 1.105 ;
      RECT 78.355 0.93 78.42 0.995 ;
      RECT 78.21 0.805 78.275 0.87 ;
      RECT 77.845 0.265 77.91 0.33 ;
      RECT 77.75 0.805 77.815 0.87 ;
      RECT 77.5825 0.265 77.6475 0.33 ;
      RECT 77.49 0.805 77.555 0.87 ;
      RECT 77.455 0.625 77.52 0.69 ;
      RECT 77.12 0.9775 77.185 1.0425 ;
      RECT 77.085 0.6 77.15 0.665 ;
      RECT 76.99 0.265 77.055 0.33 ;
      RECT 76.71 0.725 76.775 0.79 ;
      RECT 76.4 0.9775 76.465 1.0425 ;
      RECT 76.305 0.805 76.37 0.87 ;
      RECT 76.03 1.04 76.095 1.105 ;
      RECT 75.655 0.93 75.72 0.995 ;
      RECT 75.51 0.805 75.575 0.87 ;
      RECT 75.145 0.265 75.21 0.33 ;
      RECT 75.05 0.805 75.115 0.87 ;
      RECT 74.8825 0.265 74.9475 0.33 ;
      RECT 74.79 0.805 74.855 0.87 ;
      RECT 74.755 0.625 74.82 0.69 ;
      RECT 74.42 0.9775 74.485 1.0425 ;
      RECT 74.385 0.6 74.45 0.665 ;
      RECT 74.29 0.265 74.355 0.33 ;
      RECT 74.01 0.725 74.075 0.79 ;
      RECT 73.7 0.9775 73.765 1.0425 ;
      RECT 73.605 0.805 73.67 0.87 ;
      RECT 73.33 1.04 73.395 1.105 ;
      RECT 72.955 0.93 73.02 0.995 ;
      RECT 72.81 0.805 72.875 0.87 ;
      RECT 72.445 0.265 72.51 0.33 ;
      RECT 72.35 0.805 72.415 0.87 ;
      RECT 72.1825 0.265 72.2475 0.33 ;
      RECT 72.09 0.805 72.155 0.87 ;
      RECT 72.055 0.625 72.12 0.69 ;
      RECT 71.72 0.9775 71.785 1.0425 ;
      RECT 71.685 0.6 71.75 0.665 ;
      RECT 71.59 0.265 71.655 0.33 ;
      RECT 71.31 0.725 71.375 0.79 ;
      RECT 71 0.9775 71.065 1.0425 ;
      RECT 70.905 0.805 70.97 0.87 ;
      RECT 70.63 1.04 70.695 1.105 ;
      RECT 70.255 0.93 70.32 0.995 ;
      RECT 70.11 0.805 70.175 0.87 ;
      RECT 69.745 0.265 69.81 0.33 ;
      RECT 69.65 0.805 69.715 0.87 ;
      RECT 69.4825 0.265 69.5475 0.33 ;
      RECT 69.39 0.805 69.455 0.87 ;
      RECT 69.355 0.625 69.42 0.69 ;
      RECT 69.02 0.9775 69.085 1.0425 ;
      RECT 68.985 0.6 69.05 0.665 ;
      RECT 68.89 0.265 68.955 0.33 ;
      RECT 68.61 0.725 68.675 0.79 ;
      RECT 68.3 0.9775 68.365 1.0425 ;
      RECT 68.205 0.805 68.27 0.87 ;
      RECT 67.93 1.04 67.995 1.105 ;
      RECT 67.555 0.93 67.62 0.995 ;
      RECT 67.41 0.805 67.475 0.87 ;
      RECT 67.045 0.265 67.11 0.33 ;
      RECT 66.95 0.805 67.015 0.87 ;
      RECT 66.7825 0.265 66.8475 0.33 ;
      RECT 66.69 0.805 66.755 0.87 ;
      RECT 66.655 0.625 66.72 0.69 ;
      RECT 66.32 0.9775 66.385 1.0425 ;
      RECT 66.285 0.6 66.35 0.665 ;
      RECT 66.19 0.265 66.255 0.33 ;
      RECT 65.91 0.725 65.975 0.79 ;
      RECT 65.6 0.9775 65.665 1.0425 ;
      RECT 65.505 0.805 65.57 0.87 ;
      RECT 65.23 1.04 65.295 1.105 ;
      RECT 64.855 0.93 64.92 0.995 ;
      RECT 64.71 0.805 64.775 0.87 ;
      RECT 64.345 0.265 64.41 0.33 ;
      RECT 64.25 0.805 64.315 0.87 ;
      RECT 64.0825 0.265 64.1475 0.33 ;
      RECT 63.99 0.805 64.055 0.87 ;
      RECT 63.955 0.625 64.02 0.69 ;
      RECT 63.62 0.9775 63.685 1.0425 ;
      RECT 63.585 0.6 63.65 0.665 ;
      RECT 63.49 0.265 63.555 0.33 ;
      RECT 63.21 0.725 63.275 0.79 ;
      RECT 62.9 0.9775 62.965 1.0425 ;
      RECT 62.805 0.805 62.87 0.87 ;
      RECT 62.53 1.04 62.595 1.105 ;
      RECT 62.155 0.93 62.22 0.995 ;
      RECT 62.01 0.805 62.075 0.87 ;
      RECT 61.645 0.265 61.71 0.33 ;
      RECT 61.55 0.805 61.615 0.87 ;
      RECT 61.3825 0.265 61.4475 0.33 ;
      RECT 61.29 0.805 61.355 0.87 ;
      RECT 61.255 0.625 61.32 0.69 ;
      RECT 60.92 0.9775 60.985 1.0425 ;
      RECT 60.885 0.6 60.95 0.665 ;
      RECT 60.79 0.265 60.855 0.33 ;
      RECT 60.51 0.725 60.575 0.79 ;
      RECT 60.2 0.9775 60.265 1.0425 ;
      RECT 60.105 0.805 60.17 0.87 ;
      RECT 59.83 1.04 59.895 1.105 ;
      RECT 59.455 0.93 59.52 0.995 ;
      RECT 59.31 0.805 59.375 0.87 ;
      RECT 58.945 0.265 59.01 0.33 ;
      RECT 58.85 0.805 58.915 0.87 ;
      RECT 58.6825 0.265 58.7475 0.33 ;
      RECT 58.59 0.805 58.655 0.87 ;
      RECT 58.555 0.625 58.62 0.69 ;
      RECT 58.22 0.9775 58.285 1.0425 ;
      RECT 58.185 0.6 58.25 0.665 ;
      RECT 58.09 0.265 58.155 0.33 ;
      RECT 57.81 0.725 57.875 0.79 ;
      RECT 57.5 0.9775 57.565 1.0425 ;
      RECT 57.405 0.805 57.47 0.87 ;
      RECT 57.13 1.04 57.195 1.105 ;
      RECT 56.755 0.93 56.82 0.995 ;
      RECT 56.61 0.805 56.675 0.87 ;
      RECT 56.245 0.265 56.31 0.33 ;
      RECT 56.15 0.805 56.215 0.87 ;
      RECT 55.9825 0.265 56.0475 0.33 ;
      RECT 55.89 0.805 55.955 0.87 ;
      RECT 55.855 0.625 55.92 0.69 ;
      RECT 55.52 0.9775 55.585 1.0425 ;
      RECT 55.485 0.6 55.55 0.665 ;
      RECT 55.39 0.265 55.455 0.33 ;
      RECT 55.11 0.725 55.175 0.79 ;
      RECT 54.8 0.9775 54.865 1.0425 ;
      RECT 54.705 0.805 54.77 0.87 ;
      RECT 54.43 1.04 54.495 1.105 ;
      RECT 54.055 0.93 54.12 0.995 ;
      RECT 53.91 0.805 53.975 0.87 ;
      RECT 53.545 0.265 53.61 0.33 ;
      RECT 53.45 0.805 53.515 0.87 ;
      RECT 53.2825 0.265 53.3475 0.33 ;
      RECT 53.19 0.805 53.255 0.87 ;
      RECT 53.155 0.625 53.22 0.69 ;
      RECT 52.82 0.9775 52.885 1.0425 ;
      RECT 52.785 0.6 52.85 0.665 ;
      RECT 52.69 0.265 52.755 0.33 ;
      RECT 52.41 0.725 52.475 0.79 ;
      RECT 52.1 0.9775 52.165 1.0425 ;
      RECT 52.005 0.805 52.07 0.87 ;
      RECT 51.73 1.04 51.795 1.105 ;
      RECT 51.355 0.93 51.42 0.995 ;
      RECT 51.21 0.805 51.275 0.87 ;
      RECT 50.845 0.265 50.91 0.33 ;
      RECT 50.75 0.805 50.815 0.87 ;
      RECT 50.5825 0.265 50.6475 0.33 ;
      RECT 50.49 0.805 50.555 0.87 ;
      RECT 50.455 0.625 50.52 0.69 ;
      RECT 50.12 0.9775 50.185 1.0425 ;
      RECT 50.085 0.6 50.15 0.665 ;
      RECT 49.99 0.265 50.055 0.33 ;
      RECT 49.71 0.725 49.775 0.79 ;
      RECT 49.4 0.9775 49.465 1.0425 ;
      RECT 49.305 0.805 49.37 0.87 ;
      RECT 49.03 1.04 49.095 1.105 ;
      RECT 48.655 0.93 48.72 0.995 ;
      RECT 48.51 0.805 48.575 0.87 ;
      RECT 48.145 0.265 48.21 0.33 ;
      RECT 48.05 0.805 48.115 0.87 ;
      RECT 47.8825 0.265 47.9475 0.33 ;
      RECT 47.79 0.805 47.855 0.87 ;
      RECT 47.755 0.625 47.82 0.69 ;
      RECT 47.42 0.9775 47.485 1.0425 ;
      RECT 47.385 0.6 47.45 0.665 ;
      RECT 47.29 0.265 47.355 0.33 ;
      RECT 47.01 0.725 47.075 0.79 ;
      RECT 46.7 0.9775 46.765 1.0425 ;
      RECT 46.605 0.805 46.67 0.87 ;
      RECT 46.33 1.04 46.395 1.105 ;
      RECT 45.955 0.93 46.02 0.995 ;
      RECT 45.81 0.805 45.875 0.87 ;
      RECT 45.445 0.265 45.51 0.33 ;
      RECT 45.35 0.805 45.415 0.87 ;
      RECT 45.1825 0.265 45.2475 0.33 ;
      RECT 45.09 0.805 45.155 0.87 ;
      RECT 45.055 0.625 45.12 0.69 ;
      RECT 44.72 0.9775 44.785 1.0425 ;
      RECT 44.685 0.6 44.75 0.665 ;
      RECT 44.59 0.265 44.655 0.33 ;
      RECT 44.31 0.725 44.375 0.79 ;
      RECT 44 0.9775 44.065 1.0425 ;
      RECT 43.905 0.805 43.97 0.87 ;
      RECT 43.63 1.04 43.695 1.105 ;
      RECT 43.255 0.93 43.32 0.995 ;
      RECT 43.11 0.805 43.175 0.87 ;
      RECT 42.745 0.265 42.81 0.33 ;
      RECT 42.65 0.805 42.715 0.87 ;
      RECT 42.4825 0.265 42.5475 0.33 ;
      RECT 42.39 0.805 42.455 0.87 ;
      RECT 42.355 0.625 42.42 0.69 ;
      RECT 42.02 0.9775 42.085 1.0425 ;
      RECT 41.985 0.6 42.05 0.665 ;
      RECT 41.89 0.265 41.955 0.33 ;
      RECT 41.61 0.725 41.675 0.79 ;
      RECT 41.3 0.9775 41.365 1.0425 ;
      RECT 41.205 0.805 41.27 0.87 ;
      RECT 40.93 1.04 40.995 1.105 ;
      RECT 40.555 0.93 40.62 0.995 ;
      RECT 40.41 0.805 40.475 0.87 ;
      RECT 40.045 0.265 40.11 0.33 ;
      RECT 39.95 0.805 40.015 0.87 ;
      RECT 39.7825 0.265 39.8475 0.33 ;
      RECT 39.69 0.805 39.755 0.87 ;
      RECT 39.655 0.625 39.72 0.69 ;
      RECT 39.32 0.9775 39.385 1.0425 ;
      RECT 39.285 0.6 39.35 0.665 ;
      RECT 39.19 0.265 39.255 0.33 ;
      RECT 38.91 0.725 38.975 0.79 ;
      RECT 38.6 0.9775 38.665 1.0425 ;
      RECT 38.505 0.805 38.57 0.87 ;
      RECT 38.23 1.04 38.295 1.105 ;
      RECT 37.855 0.93 37.92 0.995 ;
      RECT 37.71 0.805 37.775 0.87 ;
      RECT 37.345 0.265 37.41 0.33 ;
      RECT 37.25 0.805 37.315 0.87 ;
      RECT 37.0825 0.265 37.1475 0.33 ;
      RECT 36.99 0.805 37.055 0.87 ;
      RECT 36.955 0.625 37.02 0.69 ;
      RECT 36.62 0.9775 36.685 1.0425 ;
      RECT 36.585 0.6 36.65 0.665 ;
      RECT 36.49 0.265 36.555 0.33 ;
      RECT 36.21 0.725 36.275 0.79 ;
      RECT 35.9 0.9775 35.965 1.0425 ;
      RECT 35.805 0.805 35.87 0.87 ;
      RECT 35.53 1.04 35.595 1.105 ;
      RECT 35.155 0.93 35.22 0.995 ;
      RECT 35.01 0.805 35.075 0.87 ;
      RECT 34.645 0.265 34.71 0.33 ;
      RECT 34.55 0.805 34.615 0.87 ;
      RECT 34.3825 0.265 34.4475 0.33 ;
      RECT 34.29 0.805 34.355 0.87 ;
      RECT 34.255 0.625 34.32 0.69 ;
      RECT 33.92 0.9775 33.985 1.0425 ;
      RECT 33.885 0.6 33.95 0.665 ;
      RECT 33.79 0.265 33.855 0.33 ;
      RECT 33.51 0.725 33.575 0.79 ;
      RECT 33.2 0.9775 33.265 1.0425 ;
      RECT 33.105 0.805 33.17 0.87 ;
      RECT 32.83 1.04 32.895 1.105 ;
      RECT 32.455 0.93 32.52 0.995 ;
      RECT 32.31 0.805 32.375 0.87 ;
      RECT 31.945 0.265 32.01 0.33 ;
      RECT 31.85 0.805 31.915 0.87 ;
      RECT 31.6825 0.265 31.7475 0.33 ;
      RECT 31.59 0.805 31.655 0.87 ;
      RECT 31.555 0.625 31.62 0.69 ;
      RECT 31.22 0.9775 31.285 1.0425 ;
      RECT 31.185 0.6 31.25 0.665 ;
      RECT 31.09 0.265 31.155 0.33 ;
      RECT 30.81 0.725 30.875 0.79 ;
      RECT 30.5 0.9775 30.565 1.0425 ;
      RECT 30.405 0.805 30.47 0.87 ;
      RECT 30.13 1.04 30.195 1.105 ;
      RECT 29.755 0.93 29.82 0.995 ;
      RECT 29.61 0.805 29.675 0.87 ;
      RECT 29.245 0.265 29.31 0.33 ;
      RECT 29.15 0.805 29.215 0.87 ;
      RECT 28.9825 0.265 29.0475 0.33 ;
      RECT 28.89 0.805 28.955 0.87 ;
      RECT 28.855 0.625 28.92 0.69 ;
      RECT 28.52 0.9775 28.585 1.0425 ;
      RECT 28.485 0.6 28.55 0.665 ;
      RECT 28.39 0.265 28.455 0.33 ;
      RECT 28.11 0.725 28.175 0.79 ;
      RECT 27.8 0.9775 27.865 1.0425 ;
      RECT 27.705 0.805 27.77 0.87 ;
      RECT 27.43 1.04 27.495 1.105 ;
      RECT 27.055 0.93 27.12 0.995 ;
      RECT 26.91 0.805 26.975 0.87 ;
      RECT 26.545 0.265 26.61 0.33 ;
      RECT 26.45 0.805 26.515 0.87 ;
      RECT 26.2825 0.265 26.3475 0.33 ;
      RECT 26.19 0.805 26.255 0.87 ;
      RECT 26.155 0.625 26.22 0.69 ;
      RECT 25.82 0.9775 25.885 1.0425 ;
      RECT 25.785 0.6 25.85 0.665 ;
      RECT 25.69 0.265 25.755 0.33 ;
      RECT 25.41 0.725 25.475 0.79 ;
      RECT 25.1 0.9775 25.165 1.0425 ;
      RECT 25.005 0.805 25.07 0.87 ;
      RECT 24.73 1.04 24.795 1.105 ;
      RECT 24.355 0.93 24.42 0.995 ;
      RECT 24.21 0.805 24.275 0.87 ;
      RECT 23.845 0.265 23.91 0.33 ;
      RECT 23.75 0.805 23.815 0.87 ;
      RECT 23.5825 0.265 23.6475 0.33 ;
      RECT 23.49 0.805 23.555 0.87 ;
      RECT 23.455 0.625 23.52 0.69 ;
      RECT 23.12 0.9775 23.185 1.0425 ;
      RECT 23.085 0.6 23.15 0.665 ;
      RECT 22.99 0.265 23.055 0.33 ;
      RECT 22.71 0.725 22.775 0.79 ;
      RECT 22.4 0.9775 22.465 1.0425 ;
      RECT 22.305 0.805 22.37 0.87 ;
      RECT 22.03 1.04 22.095 1.105 ;
      RECT 21.655 0.93 21.72 0.995 ;
      RECT 21.51 0.805 21.575 0.87 ;
      RECT 21.145 0.265 21.21 0.33 ;
      RECT 21.05 0.805 21.115 0.87 ;
      RECT 20.8825 0.265 20.9475 0.33 ;
      RECT 20.79 0.805 20.855 0.87 ;
      RECT 20.755 0.625 20.82 0.69 ;
      RECT 20.42 0.9775 20.485 1.0425 ;
      RECT 20.385 0.6 20.45 0.665 ;
      RECT 20.29 0.265 20.355 0.33 ;
      RECT 20.01 0.725 20.075 0.79 ;
      RECT 19.7 0.9775 19.765 1.0425 ;
      RECT 19.605 0.805 19.67 0.87 ;
      RECT 19.33 1.04 19.395 1.105 ;
      RECT 18.955 0.93 19.02 0.995 ;
      RECT 18.81 0.805 18.875 0.87 ;
      RECT 18.445 0.265 18.51 0.33 ;
      RECT 18.35 0.805 18.415 0.87 ;
      RECT 18.1825 0.265 18.2475 0.33 ;
      RECT 18.09 0.805 18.155 0.87 ;
      RECT 18.055 0.625 18.12 0.69 ;
      RECT 17.72 0.9775 17.785 1.0425 ;
      RECT 17.685 0.6 17.75 0.665 ;
      RECT 17.59 0.265 17.655 0.33 ;
      RECT 17.31 0.725 17.375 0.79 ;
      RECT 17 0.9775 17.065 1.0425 ;
      RECT 16.905 0.805 16.97 0.87 ;
      RECT 16.63 1.04 16.695 1.105 ;
      RECT 16.255 0.93 16.32 0.995 ;
      RECT 16.11 0.805 16.175 0.87 ;
      RECT 15.745 0.265 15.81 0.33 ;
      RECT 15.65 0.805 15.715 0.87 ;
      RECT 15.4825 0.265 15.5475 0.33 ;
      RECT 15.39 0.805 15.455 0.87 ;
      RECT 15.355 0.625 15.42 0.69 ;
      RECT 15.02 0.9775 15.085 1.0425 ;
      RECT 14.985 0.6 15.05 0.665 ;
      RECT 14.89 0.265 14.955 0.33 ;
      RECT 14.61 0.725 14.675 0.79 ;
      RECT 14.3 0.9775 14.365 1.0425 ;
      RECT 14.205 0.805 14.27 0.87 ;
      RECT 13.93 1.04 13.995 1.105 ;
      RECT 13.555 0.93 13.62 0.995 ;
      RECT 13.41 0.805 13.475 0.87 ;
      RECT 13.045 0.265 13.11 0.33 ;
      RECT 12.95 0.805 13.015 0.87 ;
      RECT 12.7825 0.265 12.8475 0.33 ;
      RECT 12.69 0.805 12.755 0.87 ;
      RECT 12.655 0.625 12.72 0.69 ;
      RECT 12.32 0.9775 12.385 1.0425 ;
      RECT 12.285 0.6 12.35 0.665 ;
      RECT 12.19 0.265 12.255 0.33 ;
      RECT 11.91 0.725 11.975 0.79 ;
      RECT 11.6 0.9775 11.665 1.0425 ;
      RECT 11.505 0.805 11.57 0.87 ;
      RECT 11.23 1.04 11.295 1.105 ;
      RECT 10.855 0.93 10.92 0.995 ;
      RECT 10.71 0.805 10.775 0.87 ;
      RECT 10.345 0.265 10.41 0.33 ;
      RECT 10.25 0.805 10.315 0.87 ;
      RECT 10.0825 0.265 10.1475 0.33 ;
      RECT 9.99 0.805 10.055 0.87 ;
      RECT 9.955 0.625 10.02 0.69 ;
      RECT 9.62 0.9775 9.685 1.0425 ;
      RECT 9.585 0.6 9.65 0.665 ;
      RECT 9.49 0.265 9.555 0.33 ;
      RECT 9.21 0.725 9.275 0.79 ;
      RECT 8.9 0.9775 8.965 1.0425 ;
      RECT 8.805 0.805 8.87 0.87 ;
      RECT 8.53 1.04 8.595 1.105 ;
      RECT 8.155 0.93 8.22 0.995 ;
      RECT 8.01 0.805 8.075 0.87 ;
      RECT 7.645 0.265 7.71 0.33 ;
      RECT 7.55 0.805 7.615 0.87 ;
      RECT 7.3825 0.265 7.4475 0.33 ;
      RECT 7.29 0.805 7.355 0.87 ;
      RECT 7.255 0.625 7.32 0.69 ;
      RECT 6.92 0.9775 6.985 1.0425 ;
      RECT 6.885 0.6 6.95 0.665 ;
      RECT 6.79 0.265 6.855 0.33 ;
      RECT 6.51 0.725 6.575 0.79 ;
      RECT 6.2 0.9775 6.265 1.0425 ;
      RECT 6.105 0.805 6.17 0.87 ;
      RECT 5.83 1.04 5.895 1.105 ;
      RECT 5.455 0.93 5.52 0.995 ;
      RECT 5.31 0.805 5.375 0.87 ;
      RECT 4.945 0.265 5.01 0.33 ;
      RECT 4.85 0.805 4.915 0.87 ;
      RECT 4.6825 0.265 4.7475 0.33 ;
      RECT 4.59 0.805 4.655 0.87 ;
      RECT 4.555 0.625 4.62 0.69 ;
      RECT 4.22 0.9775 4.285 1.0425 ;
      RECT 4.185 0.6 4.25 0.665 ;
      RECT 4.09 0.265 4.155 0.33 ;
      RECT 3.81 0.725 3.875 0.79 ;
      RECT 3.5 0.9775 3.565 1.0425 ;
      RECT 3.405 0.805 3.47 0.87 ;
      RECT 3.13 1.04 3.195 1.105 ;
      RECT 2.755 0.93 2.82 0.995 ;
      RECT 2.61 0.805 2.675 0.87 ;
      RECT 2.245 0.265 2.31 0.33 ;
      RECT 2.15 0.805 2.215 0.87 ;
      RECT 1.9825 0.265 2.0475 0.33 ;
      RECT 1.89 0.805 1.955 0.87 ;
      RECT 1.855 0.625 1.92 0.69 ;
      RECT 1.52 0.9775 1.585 1.0425 ;
      RECT 1.485 0.6 1.55 0.665 ;
      RECT 1.39 0.265 1.455 0.33 ;
      RECT 1.11 0.725 1.175 0.79 ;
      RECT 0.8 0.9775 0.865 1.0425 ;
      RECT 0.705 0.805 0.77 0.87 ;
      RECT 0.43 1.04 0.495 1.105 ;
      RECT 0.055 0.93 0.12 0.995 ;
    LAYER via2 ;
      RECT 87.4775 0.6225 87.5475 0.6925 ;
      RECT 85.48 0.6225 85.55 0.6925 ;
      RECT 84.7575 0.255 84.8275 0.325 ;
      RECT 84.365 0.6225 84.435 0.6925 ;
      RECT 83.2425 0.255 83.3125 0.325 ;
      RECT 82.8525 0.6225 82.9225 0.6925 ;
      RECT 80.5425 0.255 80.6125 0.325 ;
      RECT 80.1525 0.6225 80.2225 0.6925 ;
      RECT 77.8425 0.255 77.9125 0.325 ;
      RECT 77.4525 0.6225 77.5225 0.6925 ;
      RECT 75.1425 0.255 75.2125 0.325 ;
      RECT 74.7525 0.6225 74.8225 0.6925 ;
      RECT 72.4425 0.255 72.5125 0.325 ;
      RECT 72.0525 0.6225 72.1225 0.6925 ;
      RECT 69.7425 0.255 69.8125 0.325 ;
      RECT 69.3525 0.6225 69.4225 0.6925 ;
      RECT 67.0425 0.255 67.1125 0.325 ;
      RECT 66.6525 0.6225 66.7225 0.6925 ;
      RECT 64.3425 0.255 64.4125 0.325 ;
      RECT 63.9525 0.6225 64.0225 0.6925 ;
      RECT 61.6425 0.255 61.7125 0.325 ;
      RECT 61.2525 0.6225 61.3225 0.6925 ;
      RECT 58.9425 0.255 59.0125 0.325 ;
      RECT 58.5525 0.6225 58.6225 0.6925 ;
      RECT 56.2425 0.255 56.3125 0.325 ;
      RECT 55.8525 0.6225 55.9225 0.6925 ;
      RECT 53.5425 0.255 53.6125 0.325 ;
      RECT 53.1525 0.6225 53.2225 0.6925 ;
      RECT 50.8425 0.255 50.9125 0.325 ;
      RECT 50.4525 0.6225 50.5225 0.6925 ;
      RECT 48.1425 0.255 48.2125 0.325 ;
      RECT 47.7525 0.6225 47.8225 0.6925 ;
      RECT 45.4425 0.255 45.5125 0.325 ;
      RECT 45.0525 0.6225 45.1225 0.6925 ;
      RECT 42.7425 0.255 42.8125 0.325 ;
      RECT 42.3525 0.6225 42.4225 0.6925 ;
      RECT 40.0425 0.255 40.1125 0.325 ;
      RECT 39.6525 0.6225 39.7225 0.6925 ;
      RECT 37.3425 0.255 37.4125 0.325 ;
      RECT 36.9525 0.6225 37.0225 0.6925 ;
      RECT 34.6425 0.255 34.7125 0.325 ;
      RECT 34.2525 0.6225 34.3225 0.6925 ;
      RECT 31.9425 0.255 32.0125 0.325 ;
      RECT 31.5525 0.6225 31.6225 0.6925 ;
      RECT 29.2425 0.255 29.3125 0.325 ;
      RECT 28.8525 0.6225 28.9225 0.6925 ;
      RECT 26.5425 0.255 26.6125 0.325 ;
      RECT 26.1525 0.6225 26.2225 0.6925 ;
      RECT 23.8425 0.255 23.9125 0.325 ;
      RECT 23.4525 0.6225 23.5225 0.6925 ;
      RECT 21.1425 0.255 21.2125 0.325 ;
      RECT 20.7525 0.6225 20.8225 0.6925 ;
      RECT 18.4425 0.255 18.5125 0.325 ;
      RECT 18.0525 0.6225 18.1225 0.6925 ;
      RECT 15.7425 0.255 15.8125 0.325 ;
      RECT 15.3525 0.6225 15.4225 0.6925 ;
      RECT 13.0425 0.255 13.1125 0.325 ;
      RECT 12.6525 0.6225 12.7225 0.6925 ;
      RECT 10.3425 0.255 10.4125 0.325 ;
      RECT 9.9525 0.6225 10.0225 0.6925 ;
      RECT 7.6425 0.255 7.7125 0.325 ;
      RECT 7.2525 0.6225 7.3225 0.6925 ;
      RECT 4.9425 0.255 5.0125 0.325 ;
      RECT 4.5525 0.6225 4.6225 0.6925 ;
      RECT 2.2425 0.255 2.3125 0.325 ;
      RECT 1.8525 0.6225 1.9225 0.6925 ;
  END
END regfile

END LIBRARY
