* SPICE NETLIST
***************************************

.SUBCKT bit2 W R1 R2 A Z1 Z2 vss! vdd!
** N=14 EP=8 IP=0 FDC=18
M0 vss! W 1 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 4 R1 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=690 $Y=600 $D=1
M2 5 W A vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=1425 $Y=600 $D=1
M3 vss! 5 10 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=2160 $Y=600 $D=1
M4 6 10 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=2540 $Y=600 $D=1
M5 5 1 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=2985 $Y=600 $D=1
M6 6 R1 Z1 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.89e-14 AS=1.2375e-14 PD=6e-07 PS=4.55e-07 $X=3795 $Y=600 $D=1
M7 Z2 R2 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.89e-14 PD=4.55e-07 PS=6e-07 $X=4315 $Y=600 $D=1
M8 8 R2 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=5050 $Y=600 $D=1
M9 vdd! W 1 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M10 4 R1 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=690 $Y=1850 $D=0
M11 5 1 A vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=1425 $Y=1850 $D=0
M12 vdd! 5 10 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=2160 $Y=1850 $D=0
M13 6 10 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=2540 $Y=1850 $D=0
M14 5 W 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=2985 $Y=1850 $D=0
M15 6 4 Z1 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.78e-14 AS=2.475e-14 PD=7.8e-07 PS=6.35e-07 $X=3795 $Y=1850 $D=0
M16 Z2 8 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.78e-14 PD=6.35e-07 PS=7.8e-07 $X=4315 $Y=1850 $D=0
M17 8 R2 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=5050 $Y=1850 $D=0
.ENDS
***************************************
