// Global nets module 

`celldefine
module cds_globals;


supply1 vdd_;

wire vss_;


endmodule
`endcelldefine
