// Global nets module 

`celldefine
module cds_globals;


wire vss_;

supply1 vdd_;


endmodule
`endcelldefine
