* SPICE NETLIST
***************************************

.SUBCKT dff Qb CLK D Q vss! vdd!
** N=14 EP=6 IP=0 FDC=24
M0 1 CLK vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 2 1 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=970 $Y=600 $D=1
M2 9 D vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=1630 $Y=600 $D=1
M3 3 1 9 vss! NMOS_VTL L=5e-08 W=9e-08 AD=2.79e-14 AS=1.5525e-14 PD=8e-07 PS=5.25e-07 $X=2075 $Y=600 $D=1
M4 4 3 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=3155 $Y=600 $D=1
M5 10 4 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.8675e-14 AS=9e-15 PD=5.95e-07 PS=3.8e-07 $X=3815 $Y=600 $D=1
M6 3 2 10 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.8675e-14 PD=5.25e-07 PS=5.95e-07 $X=4330 $Y=600 $D=1
M7 5 2 4 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.5525e-14 PD=5.25e-07 PS=5.25e-07 $X=5280 $Y=600 $D=1
M8 Qb 5 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=6090 $Y=600 $D=1
M9 Q Qb vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=9e-15 PD=3.8e-07 PS=3.8e-07 $X=6750 $Y=600 $D=1
M10 14 Qb vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=7410 $Y=600 $D=1
M11 5 1 14 vss! NMOS_VTL L=5e-08 W=9e-08 AD=2.79e-14 AS=1.5525e-14 PD=8e-07 PS=5.25e-07 $X=7855 $Y=600 $D=1
M12 1 CLK vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=310 $Y=2055 $D=0
M13 2 1 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=970 $Y=2055 $D=0
M14 9 D vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=6.21e-14 AS=1.8e-14 PD=1.05e-06 PS=5.6e-07 $X=1630 $Y=2055 $D=0
M15 3 2 9 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=6.21e-14 PD=6.35e-07 PS=1.05e-06 $X=2420 $Y=2055 $D=0
M16 4 3 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=3155 $Y=2055 $D=0
M17 10 4 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.735e-14 AS=1.8e-14 PD=7.75e-07 PS=5.6e-07 $X=3815 $Y=2055 $D=0
M18 3 1 10 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.735e-14 PD=7.05e-07 PS=7.75e-07 $X=4330 $Y=2055 $D=0
M19 5 1 4 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=3.105e-14 PD=7.05e-07 PS=7.05e-07 $X=5280 $Y=2055 $D=0
M20 Qb 5 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=6090 $Y=2055 $D=0
M21 Q Qb vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=1.8e-14 PD=5.6e-07 PS=5.6e-07 $X=6750 $Y=2055 $D=0
M22 14 Qb vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=6.21e-14 AS=1.8e-14 PD=1.05e-06 PS=5.6e-07 $X=7410 $Y=2055 $D=0
M23 5 2 14 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=6.21e-14 PD=6.35e-07 PS=1.05e-06 $X=8200 $Y=2055 $D=0
.ENDS
***************************************
