module top_tb;

    timeunit 1ns;
    timeprecision 1ns;

    bit clk;
    always #1 clk = ~clk;

    bit rst;

            logic   [31:0]  imem_addr;
            logic   [31:0]  imem_rdata;
            logic   [31:0]  dmem_addr;
            logic           dmem_write;
            logic   [3:0]   dmem_wmask;
            logic   [31:0]  dmem_rdata;
            logic   [31:0]  dmem_wdata;

    cpu dut(.*);
    magic_dual_port mem(.*);

    mon_itf mon_itf(.*);
    monitor monitor(.itf(mon_itf));

    logic [31:0] rs1_rdata;
    logic [31:0] rd_wdata;
    logic [31:0] pc_wdata;

    // Netlist Datapath Code
    always_comb begin
        rs1_rdata[0] = dut.datapath.I0.cmp_src_a;
        rs1_rdata[1] = dut.datapath.I1.cmp_src_a;
        rs1_rdata[2] = dut.datapath.I2.cmp_src_a;
        rs1_rdata[3] = dut.datapath.I3.cmp_src_a;
        rs1_rdata[4] = dut.datapath.I4.cmp_src_a;
        rs1_rdata[5] = dut.datapath.I5.cmp_src_a;
        rs1_rdata[6] = dut.datapath.I6.cmp_src_a;
        rs1_rdata[7] = dut.datapath.I7.cmp_src_a;
        rs1_rdata[8] = dut.datapath.I8.cmp_src_a;
        rs1_rdata[9] = dut.datapath.I9.cmp_src_a;
        rs1_rdata[10] = dut.datapath.I10.cmp_src_a;
        rs1_rdata[11] = dut.datapath.I11.cmp_src_a;
        rs1_rdata[12] = dut.datapath.I12.cmp_src_a;
        rs1_rdata[13] = dut.datapath.I13.cmp_src_a;
        rs1_rdata[14] = dut.datapath.I14.cmp_src_a;
        rs1_rdata[15] = dut.datapath.I15.cmp_src_a;
        rs1_rdata[16] = dut.datapath.I16.cmp_src_a;
        rs1_rdata[17] = dut.datapath.I17.cmp_src_a;
        rs1_rdata[18] = dut.datapath.I18.cmp_src_a;
        rs1_rdata[19] = dut.datapath.I19.cmp_src_a;
        rs1_rdata[20] = dut.datapath.I20.cmp_src_a;
        rs1_rdata[21] = dut.datapath.I21.cmp_src_a;
        rs1_rdata[22] = dut.datapath.I22.cmp_src_a;
        rs1_rdata[23] = dut.datapath.I23.cmp_src_a;
        rs1_rdata[24] = dut.datapath.I24.cmp_src_a;
        rs1_rdata[25] = dut.datapath.I25.cmp_src_a;
        rs1_rdata[26] = dut.datapath.I26.cmp_src_a;
        rs1_rdata[27] = dut.datapath.I27.cmp_src_a;
        rs1_rdata[28] = dut.datapath.I28.cmp_src_a;
        rs1_rdata[29] = dut.datapath.I29.cmp_src_a;
        rs1_rdata[30] = dut.datapath.I30.cmp_src_a;
        rs1_rdata[31] = dut.datapath.I31.cmp_src_a;

        rd_wdata[0] = dut.datapath.I0.rd_mux_out;
        rd_wdata[1] = dut.datapath.I1.rd_mux_out;
        rd_wdata[2] = dut.datapath.I2.rd_mux_out;
        rd_wdata[3] = dut.datapath.I3.rd_mux_out;
        rd_wdata[4] = dut.datapath.I4.rd_mux_out;
        rd_wdata[5] = dut.datapath.I5.rd_mux_out;
        rd_wdata[6] = dut.datapath.I6.rd_mux_out;
        rd_wdata[7] = dut.datapath.I7.rd_mux_out;
        rd_wdata[8] = dut.datapath.I8.rd_mux_out;
        rd_wdata[9] = dut.datapath.I9.rd_mux_out;
        rd_wdata[10] = dut.datapath.I10.rd_mux_out;
        rd_wdata[11] = dut.datapath.I11.rd_mux_out;
        rd_wdata[12] = dut.datapath.I12.rd_mux_out;
        rd_wdata[13] = dut.datapath.I13.rd_mux_out;
        rd_wdata[14] = dut.datapath.I14.rd_mux_out;
        rd_wdata[15] = dut.datapath.I15.rd_mux_out;
        rd_wdata[16] = dut.datapath.I16.rd_mux_out;
        rd_wdata[17] = dut.datapath.I17.rd_mux_out;
        rd_wdata[18] = dut.datapath.I18.rd_mux_out;
        rd_wdata[19] = dut.datapath.I19.rd_mux_out;
        rd_wdata[20] = dut.datapath.I20.rd_mux_out;
        rd_wdata[21] = dut.datapath.I21.rd_mux_out;
        rd_wdata[22] = dut.datapath.I22.rd_mux_out;
        rd_wdata[23] = dut.datapath.I23.rd_mux_out;
        rd_wdata[24] = dut.datapath.I24.rd_mux_out;
        rd_wdata[25] = dut.datapath.I25.rd_mux_out;
        rd_wdata[26] = dut.datapath.I26.rd_mux_out;
        rd_wdata[27] = dut.datapath.I27.rd_mux_out;
        rd_wdata[28] = dut.datapath.I28.rd_mux_out;
        rd_wdata[29] = dut.datapath.I29.rd_mux_out;
        rd_wdata[30] = dut.datapath.I30.rd_mux_out;
        rd_wdata[31] = dut.datapath.I31.rd_mux_out;

        pc_wdata[0] = dut.datapath.I0.I7.pc_next;
        pc_wdata[1] = dut.datapath.I1.I7.pc_next;
        pc_wdata[2] = dut.datapath.I2.I7.pc_next;
        pc_wdata[3] = dut.datapath.I3.I7.pc_next;
        pc_wdata[4] = dut.datapath.I4.I7.pc_next;
        pc_wdata[5] = dut.datapath.I5.I7.pc_next;
        pc_wdata[6] = dut.datapath.I6.I7.pc_next;
        pc_wdata[7] = dut.datapath.I7.I7.pc_next;
        pc_wdata[8] = dut.datapath.I8.I7.pc_next;
        pc_wdata[9] = dut.datapath.I9.I7.pc_next;
        pc_wdata[10] = dut.datapath.I10.I7.pc_next;
        pc_wdata[11] = dut.datapath.I11.I7.pc_next;
        pc_wdata[12] = dut.datapath.I12.I7.pc_next;
        pc_wdata[13] = dut.datapath.I13.I7.pc_next;
        pc_wdata[14] = dut.datapath.I14.I7.pc_next;
        pc_wdata[15] = dut.datapath.I15.I7.pc_next;
        pc_wdata[16] = dut.datapath.I16.I7.pc_next;
        pc_wdata[17] = dut.datapath.I17.I7.pc_next;
        pc_wdata[18] = dut.datapath.I18.I7.pc_next;
        pc_wdata[19] = dut.datapath.I19.I7.pc_next;
        pc_wdata[20] = dut.datapath.I20.I7.pc_next;
        pc_wdata[21] = dut.datapath.I21.I7.pc_next;
        pc_wdata[22] = dut.datapath.I22.I7.pc_next;
        pc_wdata[23] = dut.datapath.I23.I7.pc_next;
        pc_wdata[24] = dut.datapath.I24.I7.pc_next;
        pc_wdata[25] = dut.datapath.I25.I7.pc_next;
        pc_wdata[26] = dut.datapath.I26.I7.pc_next;
        pc_wdata[27] = dut.datapath.I27.I7.pc_next;
        pc_wdata[28] = dut.datapath.I28.I7.pc_next;
        pc_wdata[29] = dut.datapath.I29.I7.pc_next;
        pc_wdata[30] = dut.datapath.I30.I7.pc_next;
        pc_wdata[31] = dut.datapath.I31.I7.pc_next;
    end

    // Netlist Datapath Code
    logic [31:0] real_rf_data[32];
    always_comb begin
        for (int j = 0; j < 32; j++) begin
            real_rf_data[0][j] = 1'b0;
        end

        real_rf_data[1][0] = dut.datapath.I0.I9.I0.I1.Bit;
        real_rf_data[1][1] = dut.datapath.I1.I9.I0.I1.Bit;
        real_rf_data[1][2] = dut.datapath.I2.I9.I0.I1.Bit;
        real_rf_data[1][3] = dut.datapath.I3.I9.I0.I1.Bit;
        real_rf_data[1][4] = dut.datapath.I4.I9.I0.I1.Bit;
        real_rf_data[1][5] = dut.datapath.I5.I9.I0.I1.Bit;
        real_rf_data[1][6] = dut.datapath.I6.I9.I0.I1.Bit;
        real_rf_data[1][7] = dut.datapath.I7.I9.I0.I1.Bit;
        real_rf_data[1][8] = dut.datapath.I8.I9.I0.I1.Bit;
        real_rf_data[1][9] = dut.datapath.I9.I9.I0.I1.Bit;
        real_rf_data[1][10] = dut.datapath.I10.I9.I0.I1.Bit;
        real_rf_data[1][11] = dut.datapath.I11.I9.I0.I1.Bit;
        real_rf_data[1][12] = dut.datapath.I12.I9.I0.I1.Bit;
        real_rf_data[1][13] = dut.datapath.I13.I9.I0.I1.Bit;
        real_rf_data[1][14] = dut.datapath.I14.I9.I0.I1.Bit;
        real_rf_data[1][15] = dut.datapath.I15.I9.I0.I1.Bit;
        real_rf_data[1][16] = dut.datapath.I16.I9.I0.I1.Bit;
        real_rf_data[1][17] = dut.datapath.I17.I9.I0.I1.Bit;
        real_rf_data[1][18] = dut.datapath.I18.I9.I0.I1.Bit;
        real_rf_data[1][19] = dut.datapath.I19.I9.I0.I1.Bit;
        real_rf_data[1][20] = dut.datapath.I20.I9.I0.I1.Bit;
        real_rf_data[1][21] = dut.datapath.I21.I9.I0.I1.Bit;
        real_rf_data[1][22] = dut.datapath.I22.I9.I0.I1.Bit;
        real_rf_data[1][23] = dut.datapath.I23.I9.I0.I1.Bit;
        real_rf_data[1][24] = dut.datapath.I24.I9.I0.I1.Bit;
        real_rf_data[1][25] = dut.datapath.I25.I9.I0.I1.Bit;
        real_rf_data[1][26] = dut.datapath.I26.I9.I0.I1.Bit;
        real_rf_data[1][27] = dut.datapath.I27.I9.I0.I1.Bit;
        real_rf_data[1][28] = dut.datapath.I28.I9.I0.I1.Bit;
        real_rf_data[1][29] = dut.datapath.I29.I9.I0.I1.Bit;
        real_rf_data[1][30] = dut.datapath.I30.I9.I0.I1.Bit;
        real_rf_data[1][31] = dut.datapath.I31.I9.I0.I1.Bit;
        real_rf_data[2][0] = dut.datapath.I0.I9.I0.I2.Bit;
        real_rf_data[2][1] = dut.datapath.I1.I9.I0.I2.Bit;
        real_rf_data[2][2] = dut.datapath.I2.I9.I0.I2.Bit;
        real_rf_data[2][3] = dut.datapath.I3.I9.I0.I2.Bit;
        real_rf_data[2][4] = dut.datapath.I4.I9.I0.I2.Bit;
        real_rf_data[2][5] = dut.datapath.I5.I9.I0.I2.Bit;
        real_rf_data[2][6] = dut.datapath.I6.I9.I0.I2.Bit;
        real_rf_data[2][7] = dut.datapath.I7.I9.I0.I2.Bit;
        real_rf_data[2][8] = dut.datapath.I8.I9.I0.I2.Bit;
        real_rf_data[2][9] = dut.datapath.I9.I9.I0.I2.Bit;
        real_rf_data[2][10] = dut.datapath.I10.I9.I0.I2.Bit;
        real_rf_data[2][11] = dut.datapath.I11.I9.I0.I2.Bit;
        real_rf_data[2][12] = dut.datapath.I12.I9.I0.I2.Bit;
        real_rf_data[2][13] = dut.datapath.I13.I9.I0.I2.Bit;
        real_rf_data[2][14] = dut.datapath.I14.I9.I0.I2.Bit;
        real_rf_data[2][15] = dut.datapath.I15.I9.I0.I2.Bit;
        real_rf_data[2][16] = dut.datapath.I16.I9.I0.I2.Bit;
        real_rf_data[2][17] = dut.datapath.I17.I9.I0.I2.Bit;
        real_rf_data[2][18] = dut.datapath.I18.I9.I0.I2.Bit;
        real_rf_data[2][19] = dut.datapath.I19.I9.I0.I2.Bit;
        real_rf_data[2][20] = dut.datapath.I20.I9.I0.I2.Bit;
        real_rf_data[2][21] = dut.datapath.I21.I9.I0.I2.Bit;
        real_rf_data[2][22] = dut.datapath.I22.I9.I0.I2.Bit;
        real_rf_data[2][23] = dut.datapath.I23.I9.I0.I2.Bit;
        real_rf_data[2][24] = dut.datapath.I24.I9.I0.I2.Bit;
        real_rf_data[2][25] = dut.datapath.I25.I9.I0.I2.Bit;
        real_rf_data[2][26] = dut.datapath.I26.I9.I0.I2.Bit;
        real_rf_data[2][27] = dut.datapath.I27.I9.I0.I2.Bit;
        real_rf_data[2][28] = dut.datapath.I28.I9.I0.I2.Bit;
        real_rf_data[2][29] = dut.datapath.I29.I9.I0.I2.Bit;
        real_rf_data[2][30] = dut.datapath.I30.I9.I0.I2.Bit;
        real_rf_data[2][31] = dut.datapath.I31.I9.I0.I2.Bit;
        real_rf_data[3][0] = dut.datapath.I0.I9.I0.I3.Bit;
        real_rf_data[3][1] = dut.datapath.I1.I9.I0.I3.Bit;
        real_rf_data[3][2] = dut.datapath.I2.I9.I0.I3.Bit;
        real_rf_data[3][3] = dut.datapath.I3.I9.I0.I3.Bit;
        real_rf_data[3][4] = dut.datapath.I4.I9.I0.I3.Bit;
        real_rf_data[3][5] = dut.datapath.I5.I9.I0.I3.Bit;
        real_rf_data[3][6] = dut.datapath.I6.I9.I0.I3.Bit;
        real_rf_data[3][7] = dut.datapath.I7.I9.I0.I3.Bit;
        real_rf_data[3][8] = dut.datapath.I8.I9.I0.I3.Bit;
        real_rf_data[3][9] = dut.datapath.I9.I9.I0.I3.Bit;
        real_rf_data[3][10] = dut.datapath.I10.I9.I0.I3.Bit;
        real_rf_data[3][11] = dut.datapath.I11.I9.I0.I3.Bit;
        real_rf_data[3][12] = dut.datapath.I12.I9.I0.I3.Bit;
        real_rf_data[3][13] = dut.datapath.I13.I9.I0.I3.Bit;
        real_rf_data[3][14] = dut.datapath.I14.I9.I0.I3.Bit;
        real_rf_data[3][15] = dut.datapath.I15.I9.I0.I3.Bit;
        real_rf_data[3][16] = dut.datapath.I16.I9.I0.I3.Bit;
        real_rf_data[3][17] = dut.datapath.I17.I9.I0.I3.Bit;
        real_rf_data[3][18] = dut.datapath.I18.I9.I0.I3.Bit;
        real_rf_data[3][19] = dut.datapath.I19.I9.I0.I3.Bit;
        real_rf_data[3][20] = dut.datapath.I20.I9.I0.I3.Bit;
        real_rf_data[3][21] = dut.datapath.I21.I9.I0.I3.Bit;
        real_rf_data[3][22] = dut.datapath.I22.I9.I0.I3.Bit;
        real_rf_data[3][23] = dut.datapath.I23.I9.I0.I3.Bit;
        real_rf_data[3][24] = dut.datapath.I24.I9.I0.I3.Bit;
        real_rf_data[3][25] = dut.datapath.I25.I9.I0.I3.Bit;
        real_rf_data[3][26] = dut.datapath.I26.I9.I0.I3.Bit;
        real_rf_data[3][27] = dut.datapath.I27.I9.I0.I3.Bit;
        real_rf_data[3][28] = dut.datapath.I28.I9.I0.I3.Bit;
        real_rf_data[3][29] = dut.datapath.I29.I9.I0.I3.Bit;
        real_rf_data[3][30] = dut.datapath.I30.I9.I0.I3.Bit;
        real_rf_data[3][31] = dut.datapath.I31.I9.I0.I3.Bit;
        real_rf_data[4][0] = dut.datapath.I0.I9.I0.I4.Bit;
        real_rf_data[4][1] = dut.datapath.I1.I9.I0.I4.Bit;
        real_rf_data[4][2] = dut.datapath.I2.I9.I0.I4.Bit;
        real_rf_data[4][3] = dut.datapath.I3.I9.I0.I4.Bit;
        real_rf_data[4][4] = dut.datapath.I4.I9.I0.I4.Bit;
        real_rf_data[4][5] = dut.datapath.I5.I9.I0.I4.Bit;
        real_rf_data[4][6] = dut.datapath.I6.I9.I0.I4.Bit;
        real_rf_data[4][7] = dut.datapath.I7.I9.I0.I4.Bit;
        real_rf_data[4][8] = dut.datapath.I8.I9.I0.I4.Bit;
        real_rf_data[4][9] = dut.datapath.I9.I9.I0.I4.Bit;
        real_rf_data[4][10] = dut.datapath.I10.I9.I0.I4.Bit;
        real_rf_data[4][11] = dut.datapath.I11.I9.I0.I4.Bit;
        real_rf_data[4][12] = dut.datapath.I12.I9.I0.I4.Bit;
        real_rf_data[4][13] = dut.datapath.I13.I9.I0.I4.Bit;
        real_rf_data[4][14] = dut.datapath.I14.I9.I0.I4.Bit;
        real_rf_data[4][15] = dut.datapath.I15.I9.I0.I4.Bit;
        real_rf_data[4][16] = dut.datapath.I16.I9.I0.I4.Bit;
        real_rf_data[4][17] = dut.datapath.I17.I9.I0.I4.Bit;
        real_rf_data[4][18] = dut.datapath.I18.I9.I0.I4.Bit;
        real_rf_data[4][19] = dut.datapath.I19.I9.I0.I4.Bit;
        real_rf_data[4][20] = dut.datapath.I20.I9.I0.I4.Bit;
        real_rf_data[4][21] = dut.datapath.I21.I9.I0.I4.Bit;
        real_rf_data[4][22] = dut.datapath.I22.I9.I0.I4.Bit;
        real_rf_data[4][23] = dut.datapath.I23.I9.I0.I4.Bit;
        real_rf_data[4][24] = dut.datapath.I24.I9.I0.I4.Bit;
        real_rf_data[4][25] = dut.datapath.I25.I9.I0.I4.Bit;
        real_rf_data[4][26] = dut.datapath.I26.I9.I0.I4.Bit;
        real_rf_data[4][27] = dut.datapath.I27.I9.I0.I4.Bit;
        real_rf_data[4][28] = dut.datapath.I28.I9.I0.I4.Bit;
        real_rf_data[4][29] = dut.datapath.I29.I9.I0.I4.Bit;
        real_rf_data[4][30] = dut.datapath.I30.I9.I0.I4.Bit;
        real_rf_data[4][31] = dut.datapath.I31.I9.I0.I4.Bit;
        real_rf_data[5][0] = dut.datapath.I0.I9.I0.I5.Bit;
        real_rf_data[5][1] = dut.datapath.I1.I9.I0.I5.Bit;
        real_rf_data[5][2] = dut.datapath.I2.I9.I0.I5.Bit;
        real_rf_data[5][3] = dut.datapath.I3.I9.I0.I5.Bit;
        real_rf_data[5][4] = dut.datapath.I4.I9.I0.I5.Bit;
        real_rf_data[5][5] = dut.datapath.I5.I9.I0.I5.Bit;
        real_rf_data[5][6] = dut.datapath.I6.I9.I0.I5.Bit;
        real_rf_data[5][7] = dut.datapath.I7.I9.I0.I5.Bit;
        real_rf_data[5][8] = dut.datapath.I8.I9.I0.I5.Bit;
        real_rf_data[5][9] = dut.datapath.I9.I9.I0.I5.Bit;
        real_rf_data[5][10] = dut.datapath.I10.I9.I0.I5.Bit;
        real_rf_data[5][11] = dut.datapath.I11.I9.I0.I5.Bit;
        real_rf_data[5][12] = dut.datapath.I12.I9.I0.I5.Bit;
        real_rf_data[5][13] = dut.datapath.I13.I9.I0.I5.Bit;
        real_rf_data[5][14] = dut.datapath.I14.I9.I0.I5.Bit;
        real_rf_data[5][15] = dut.datapath.I15.I9.I0.I5.Bit;
        real_rf_data[5][16] = dut.datapath.I16.I9.I0.I5.Bit;
        real_rf_data[5][17] = dut.datapath.I17.I9.I0.I5.Bit;
        real_rf_data[5][18] = dut.datapath.I18.I9.I0.I5.Bit;
        real_rf_data[5][19] = dut.datapath.I19.I9.I0.I5.Bit;
        real_rf_data[5][20] = dut.datapath.I20.I9.I0.I5.Bit;
        real_rf_data[5][21] = dut.datapath.I21.I9.I0.I5.Bit;
        real_rf_data[5][22] = dut.datapath.I22.I9.I0.I5.Bit;
        real_rf_data[5][23] = dut.datapath.I23.I9.I0.I5.Bit;
        real_rf_data[5][24] = dut.datapath.I24.I9.I0.I5.Bit;
        real_rf_data[5][25] = dut.datapath.I25.I9.I0.I5.Bit;
        real_rf_data[5][26] = dut.datapath.I26.I9.I0.I5.Bit;
        real_rf_data[5][27] = dut.datapath.I27.I9.I0.I5.Bit;
        real_rf_data[5][28] = dut.datapath.I28.I9.I0.I5.Bit;
        real_rf_data[5][29] = dut.datapath.I29.I9.I0.I5.Bit;
        real_rf_data[5][30] = dut.datapath.I30.I9.I0.I5.Bit;
        real_rf_data[5][31] = dut.datapath.I31.I9.I0.I5.Bit;
        real_rf_data[6][0] = dut.datapath.I0.I9.I0.I6.Bit;
        real_rf_data[6][1] = dut.datapath.I1.I9.I0.I6.Bit;
        real_rf_data[6][2] = dut.datapath.I2.I9.I0.I6.Bit;
        real_rf_data[6][3] = dut.datapath.I3.I9.I0.I6.Bit;
        real_rf_data[6][4] = dut.datapath.I4.I9.I0.I6.Bit;
        real_rf_data[6][5] = dut.datapath.I5.I9.I0.I6.Bit;
        real_rf_data[6][6] = dut.datapath.I6.I9.I0.I6.Bit;
        real_rf_data[6][7] = dut.datapath.I7.I9.I0.I6.Bit;
        real_rf_data[6][8] = dut.datapath.I8.I9.I0.I6.Bit;
        real_rf_data[6][9] = dut.datapath.I9.I9.I0.I6.Bit;
        real_rf_data[6][10] = dut.datapath.I10.I9.I0.I6.Bit;
        real_rf_data[6][11] = dut.datapath.I11.I9.I0.I6.Bit;
        real_rf_data[6][12] = dut.datapath.I12.I9.I0.I6.Bit;
        real_rf_data[6][13] = dut.datapath.I13.I9.I0.I6.Bit;
        real_rf_data[6][14] = dut.datapath.I14.I9.I0.I6.Bit;
        real_rf_data[6][15] = dut.datapath.I15.I9.I0.I6.Bit;
        real_rf_data[6][16] = dut.datapath.I16.I9.I0.I6.Bit;
        real_rf_data[6][17] = dut.datapath.I17.I9.I0.I6.Bit;
        real_rf_data[6][18] = dut.datapath.I18.I9.I0.I6.Bit;
        real_rf_data[6][19] = dut.datapath.I19.I9.I0.I6.Bit;
        real_rf_data[6][20] = dut.datapath.I20.I9.I0.I6.Bit;
        real_rf_data[6][21] = dut.datapath.I21.I9.I0.I6.Bit;
        real_rf_data[6][22] = dut.datapath.I22.I9.I0.I6.Bit;
        real_rf_data[6][23] = dut.datapath.I23.I9.I0.I6.Bit;
        real_rf_data[6][24] = dut.datapath.I24.I9.I0.I6.Bit;
        real_rf_data[6][25] = dut.datapath.I25.I9.I0.I6.Bit;
        real_rf_data[6][26] = dut.datapath.I26.I9.I0.I6.Bit;
        real_rf_data[6][27] = dut.datapath.I27.I9.I0.I6.Bit;
        real_rf_data[6][28] = dut.datapath.I28.I9.I0.I6.Bit;
        real_rf_data[6][29] = dut.datapath.I29.I9.I0.I6.Bit;
        real_rf_data[6][30] = dut.datapath.I30.I9.I0.I6.Bit;
        real_rf_data[6][31] = dut.datapath.I31.I9.I0.I6.Bit;
        real_rf_data[7][0] = dut.datapath.I0.I9.I0.I7.Bit;
        real_rf_data[7][1] = dut.datapath.I1.I9.I0.I7.Bit;
        real_rf_data[7][2] = dut.datapath.I2.I9.I0.I7.Bit;
        real_rf_data[7][3] = dut.datapath.I3.I9.I0.I7.Bit;
        real_rf_data[7][4] = dut.datapath.I4.I9.I0.I7.Bit;
        real_rf_data[7][5] = dut.datapath.I5.I9.I0.I7.Bit;
        real_rf_data[7][6] = dut.datapath.I6.I9.I0.I7.Bit;
        real_rf_data[7][7] = dut.datapath.I7.I9.I0.I7.Bit;
        real_rf_data[7][8] = dut.datapath.I8.I9.I0.I7.Bit;
        real_rf_data[7][9] = dut.datapath.I9.I9.I0.I7.Bit;
        real_rf_data[7][10] = dut.datapath.I10.I9.I0.I7.Bit;
        real_rf_data[7][11] = dut.datapath.I11.I9.I0.I7.Bit;
        real_rf_data[7][12] = dut.datapath.I12.I9.I0.I7.Bit;
        real_rf_data[7][13] = dut.datapath.I13.I9.I0.I7.Bit;
        real_rf_data[7][14] = dut.datapath.I14.I9.I0.I7.Bit;
        real_rf_data[7][15] = dut.datapath.I15.I9.I0.I7.Bit;
        real_rf_data[7][16] = dut.datapath.I16.I9.I0.I7.Bit;
        real_rf_data[7][17] = dut.datapath.I17.I9.I0.I7.Bit;
        real_rf_data[7][18] = dut.datapath.I18.I9.I0.I7.Bit;
        real_rf_data[7][19] = dut.datapath.I19.I9.I0.I7.Bit;
        real_rf_data[7][20] = dut.datapath.I20.I9.I0.I7.Bit;
        real_rf_data[7][21] = dut.datapath.I21.I9.I0.I7.Bit;
        real_rf_data[7][22] = dut.datapath.I22.I9.I0.I7.Bit;
        real_rf_data[7][23] = dut.datapath.I23.I9.I0.I7.Bit;
        real_rf_data[7][24] = dut.datapath.I24.I9.I0.I7.Bit;
        real_rf_data[7][25] = dut.datapath.I25.I9.I0.I7.Bit;
        real_rf_data[7][26] = dut.datapath.I26.I9.I0.I7.Bit;
        real_rf_data[7][27] = dut.datapath.I27.I9.I0.I7.Bit;
        real_rf_data[7][28] = dut.datapath.I28.I9.I0.I7.Bit;
        real_rf_data[7][29] = dut.datapath.I29.I9.I0.I7.Bit;
        real_rf_data[7][30] = dut.datapath.I30.I9.I0.I7.Bit;
        real_rf_data[7][31] = dut.datapath.I31.I9.I0.I7.Bit;
        real_rf_data[8][0] = dut.datapath.I0.I9.I0.I8.Bit;
        real_rf_data[8][1] = dut.datapath.I1.I9.I0.I8.Bit;
        real_rf_data[8][2] = dut.datapath.I2.I9.I0.I8.Bit;
        real_rf_data[8][3] = dut.datapath.I3.I9.I0.I8.Bit;
        real_rf_data[8][4] = dut.datapath.I4.I9.I0.I8.Bit;
        real_rf_data[8][5] = dut.datapath.I5.I9.I0.I8.Bit;
        real_rf_data[8][6] = dut.datapath.I6.I9.I0.I8.Bit;
        real_rf_data[8][7] = dut.datapath.I7.I9.I0.I8.Bit;
        real_rf_data[8][8] = dut.datapath.I8.I9.I0.I8.Bit;
        real_rf_data[8][9] = dut.datapath.I9.I9.I0.I8.Bit;
        real_rf_data[8][10] = dut.datapath.I10.I9.I0.I8.Bit;
        real_rf_data[8][11] = dut.datapath.I11.I9.I0.I8.Bit;
        real_rf_data[8][12] = dut.datapath.I12.I9.I0.I8.Bit;
        real_rf_data[8][13] = dut.datapath.I13.I9.I0.I8.Bit;
        real_rf_data[8][14] = dut.datapath.I14.I9.I0.I8.Bit;
        real_rf_data[8][15] = dut.datapath.I15.I9.I0.I8.Bit;
        real_rf_data[8][16] = dut.datapath.I16.I9.I0.I8.Bit;
        real_rf_data[8][17] = dut.datapath.I17.I9.I0.I8.Bit;
        real_rf_data[8][18] = dut.datapath.I18.I9.I0.I8.Bit;
        real_rf_data[8][19] = dut.datapath.I19.I9.I0.I8.Bit;
        real_rf_data[8][20] = dut.datapath.I20.I9.I0.I8.Bit;
        real_rf_data[8][21] = dut.datapath.I21.I9.I0.I8.Bit;
        real_rf_data[8][22] = dut.datapath.I22.I9.I0.I8.Bit;
        real_rf_data[8][23] = dut.datapath.I23.I9.I0.I8.Bit;
        real_rf_data[8][24] = dut.datapath.I24.I9.I0.I8.Bit;
        real_rf_data[8][25] = dut.datapath.I25.I9.I0.I8.Bit;
        real_rf_data[8][26] = dut.datapath.I26.I9.I0.I8.Bit;
        real_rf_data[8][27] = dut.datapath.I27.I9.I0.I8.Bit;
        real_rf_data[8][28] = dut.datapath.I28.I9.I0.I8.Bit;
        real_rf_data[8][29] = dut.datapath.I29.I9.I0.I8.Bit;
        real_rf_data[8][30] = dut.datapath.I30.I9.I0.I8.Bit;
        real_rf_data[8][31] = dut.datapath.I31.I9.I0.I8.Bit;
        real_rf_data[9][0] = dut.datapath.I0.I9.I0.I9.Bit;
        real_rf_data[9][1] = dut.datapath.I1.I9.I0.I9.Bit;
        real_rf_data[9][2] = dut.datapath.I2.I9.I0.I9.Bit;
        real_rf_data[9][3] = dut.datapath.I3.I9.I0.I9.Bit;
        real_rf_data[9][4] = dut.datapath.I4.I9.I0.I9.Bit;
        real_rf_data[9][5] = dut.datapath.I5.I9.I0.I9.Bit;
        real_rf_data[9][6] = dut.datapath.I6.I9.I0.I9.Bit;
        real_rf_data[9][7] = dut.datapath.I7.I9.I0.I9.Bit;
        real_rf_data[9][8] = dut.datapath.I8.I9.I0.I9.Bit;
        real_rf_data[9][9] = dut.datapath.I9.I9.I0.I9.Bit;
        real_rf_data[9][10] = dut.datapath.I10.I9.I0.I9.Bit;
        real_rf_data[9][11] = dut.datapath.I11.I9.I0.I9.Bit;
        real_rf_data[9][12] = dut.datapath.I12.I9.I0.I9.Bit;
        real_rf_data[9][13] = dut.datapath.I13.I9.I0.I9.Bit;
        real_rf_data[9][14] = dut.datapath.I14.I9.I0.I9.Bit;
        real_rf_data[9][15] = dut.datapath.I15.I9.I0.I9.Bit;
        real_rf_data[9][16] = dut.datapath.I16.I9.I0.I9.Bit;
        real_rf_data[9][17] = dut.datapath.I17.I9.I0.I9.Bit;
        real_rf_data[9][18] = dut.datapath.I18.I9.I0.I9.Bit;
        real_rf_data[9][19] = dut.datapath.I19.I9.I0.I9.Bit;
        real_rf_data[9][20] = dut.datapath.I20.I9.I0.I9.Bit;
        real_rf_data[9][21] = dut.datapath.I21.I9.I0.I9.Bit;
        real_rf_data[9][22] = dut.datapath.I22.I9.I0.I9.Bit;
        real_rf_data[9][23] = dut.datapath.I23.I9.I0.I9.Bit;
        real_rf_data[9][24] = dut.datapath.I24.I9.I0.I9.Bit;
        real_rf_data[9][25] = dut.datapath.I25.I9.I0.I9.Bit;
        real_rf_data[9][26] = dut.datapath.I26.I9.I0.I9.Bit;
        real_rf_data[9][27] = dut.datapath.I27.I9.I0.I9.Bit;
        real_rf_data[9][28] = dut.datapath.I28.I9.I0.I9.Bit;
        real_rf_data[9][29] = dut.datapath.I29.I9.I0.I9.Bit;
        real_rf_data[9][30] = dut.datapath.I30.I9.I0.I9.Bit;
        real_rf_data[9][31] = dut.datapath.I31.I9.I0.I9.Bit;
        real_rf_data[10][0] = dut.datapath.I0.I9.I0.I10.Bit;
        real_rf_data[10][1] = dut.datapath.I1.I9.I0.I10.Bit;
        real_rf_data[10][2] = dut.datapath.I2.I9.I0.I10.Bit;
        real_rf_data[10][3] = dut.datapath.I3.I9.I0.I10.Bit;
        real_rf_data[10][4] = dut.datapath.I4.I9.I0.I10.Bit;
        real_rf_data[10][5] = dut.datapath.I5.I9.I0.I10.Bit;
        real_rf_data[10][6] = dut.datapath.I6.I9.I0.I10.Bit;
        real_rf_data[10][7] = dut.datapath.I7.I9.I0.I10.Bit;
        real_rf_data[10][8] = dut.datapath.I8.I9.I0.I10.Bit;
        real_rf_data[10][9] = dut.datapath.I9.I9.I0.I10.Bit;
        real_rf_data[10][10] = dut.datapath.I10.I9.I0.I10.Bit;
        real_rf_data[10][11] = dut.datapath.I11.I9.I0.I10.Bit;
        real_rf_data[10][12] = dut.datapath.I12.I9.I0.I10.Bit;
        real_rf_data[10][13] = dut.datapath.I13.I9.I0.I10.Bit;
        real_rf_data[10][14] = dut.datapath.I14.I9.I0.I10.Bit;
        real_rf_data[10][15] = dut.datapath.I15.I9.I0.I10.Bit;
        real_rf_data[10][16] = dut.datapath.I16.I9.I0.I10.Bit;
        real_rf_data[10][17] = dut.datapath.I17.I9.I0.I10.Bit;
        real_rf_data[10][18] = dut.datapath.I18.I9.I0.I10.Bit;
        real_rf_data[10][19] = dut.datapath.I19.I9.I0.I10.Bit;
        real_rf_data[10][20] = dut.datapath.I20.I9.I0.I10.Bit;
        real_rf_data[10][21] = dut.datapath.I21.I9.I0.I10.Bit;
        real_rf_data[10][22] = dut.datapath.I22.I9.I0.I10.Bit;
        real_rf_data[10][23] = dut.datapath.I23.I9.I0.I10.Bit;
        real_rf_data[10][24] = dut.datapath.I24.I9.I0.I10.Bit;
        real_rf_data[10][25] = dut.datapath.I25.I9.I0.I10.Bit;
        real_rf_data[10][26] = dut.datapath.I26.I9.I0.I10.Bit;
        real_rf_data[10][27] = dut.datapath.I27.I9.I0.I10.Bit;
        real_rf_data[10][28] = dut.datapath.I28.I9.I0.I10.Bit;
        real_rf_data[10][29] = dut.datapath.I29.I9.I0.I10.Bit;
        real_rf_data[10][30] = dut.datapath.I30.I9.I0.I10.Bit;
        real_rf_data[10][31] = dut.datapath.I31.I9.I0.I10.Bit;
        real_rf_data[11][0] = dut.datapath.I0.I9.I0.I11.Bit;
        real_rf_data[11][1] = dut.datapath.I1.I9.I0.I11.Bit;
        real_rf_data[11][2] = dut.datapath.I2.I9.I0.I11.Bit;
        real_rf_data[11][3] = dut.datapath.I3.I9.I0.I11.Bit;
        real_rf_data[11][4] = dut.datapath.I4.I9.I0.I11.Bit;
        real_rf_data[11][5] = dut.datapath.I5.I9.I0.I11.Bit;
        real_rf_data[11][6] = dut.datapath.I6.I9.I0.I11.Bit;
        real_rf_data[11][7] = dut.datapath.I7.I9.I0.I11.Bit;
        real_rf_data[11][8] = dut.datapath.I8.I9.I0.I11.Bit;
        real_rf_data[11][9] = dut.datapath.I9.I9.I0.I11.Bit;
        real_rf_data[11][10] = dut.datapath.I10.I9.I0.I11.Bit;
        real_rf_data[11][11] = dut.datapath.I11.I9.I0.I11.Bit;
        real_rf_data[11][12] = dut.datapath.I12.I9.I0.I11.Bit;
        real_rf_data[11][13] = dut.datapath.I13.I9.I0.I11.Bit;
        real_rf_data[11][14] = dut.datapath.I14.I9.I0.I11.Bit;
        real_rf_data[11][15] = dut.datapath.I15.I9.I0.I11.Bit;
        real_rf_data[11][16] = dut.datapath.I16.I9.I0.I11.Bit;
        real_rf_data[11][17] = dut.datapath.I17.I9.I0.I11.Bit;
        real_rf_data[11][18] = dut.datapath.I18.I9.I0.I11.Bit;
        real_rf_data[11][19] = dut.datapath.I19.I9.I0.I11.Bit;
        real_rf_data[11][20] = dut.datapath.I20.I9.I0.I11.Bit;
        real_rf_data[11][21] = dut.datapath.I21.I9.I0.I11.Bit;
        real_rf_data[11][22] = dut.datapath.I22.I9.I0.I11.Bit;
        real_rf_data[11][23] = dut.datapath.I23.I9.I0.I11.Bit;
        real_rf_data[11][24] = dut.datapath.I24.I9.I0.I11.Bit;
        real_rf_data[11][25] = dut.datapath.I25.I9.I0.I11.Bit;
        real_rf_data[11][26] = dut.datapath.I26.I9.I0.I11.Bit;
        real_rf_data[11][27] = dut.datapath.I27.I9.I0.I11.Bit;
        real_rf_data[11][28] = dut.datapath.I28.I9.I0.I11.Bit;
        real_rf_data[11][29] = dut.datapath.I29.I9.I0.I11.Bit;
        real_rf_data[11][30] = dut.datapath.I30.I9.I0.I11.Bit;
        real_rf_data[11][31] = dut.datapath.I31.I9.I0.I11.Bit;
        real_rf_data[12][0] = dut.datapath.I0.I9.I0.I12.Bit;
        real_rf_data[12][1] = dut.datapath.I1.I9.I0.I12.Bit;
        real_rf_data[12][2] = dut.datapath.I2.I9.I0.I12.Bit;
        real_rf_data[12][3] = dut.datapath.I3.I9.I0.I12.Bit;
        real_rf_data[12][4] = dut.datapath.I4.I9.I0.I12.Bit;
        real_rf_data[12][5] = dut.datapath.I5.I9.I0.I12.Bit;
        real_rf_data[12][6] = dut.datapath.I6.I9.I0.I12.Bit;
        real_rf_data[12][7] = dut.datapath.I7.I9.I0.I12.Bit;
        real_rf_data[12][8] = dut.datapath.I8.I9.I0.I12.Bit;
        real_rf_data[12][9] = dut.datapath.I9.I9.I0.I12.Bit;
        real_rf_data[12][10] = dut.datapath.I10.I9.I0.I12.Bit;
        real_rf_data[12][11] = dut.datapath.I11.I9.I0.I12.Bit;
        real_rf_data[12][12] = dut.datapath.I12.I9.I0.I12.Bit;
        real_rf_data[12][13] = dut.datapath.I13.I9.I0.I12.Bit;
        real_rf_data[12][14] = dut.datapath.I14.I9.I0.I12.Bit;
        real_rf_data[12][15] = dut.datapath.I15.I9.I0.I12.Bit;
        real_rf_data[12][16] = dut.datapath.I16.I9.I0.I12.Bit;
        real_rf_data[12][17] = dut.datapath.I17.I9.I0.I12.Bit;
        real_rf_data[12][18] = dut.datapath.I18.I9.I0.I12.Bit;
        real_rf_data[12][19] = dut.datapath.I19.I9.I0.I12.Bit;
        real_rf_data[12][20] = dut.datapath.I20.I9.I0.I12.Bit;
        real_rf_data[12][21] = dut.datapath.I21.I9.I0.I12.Bit;
        real_rf_data[12][22] = dut.datapath.I22.I9.I0.I12.Bit;
        real_rf_data[12][23] = dut.datapath.I23.I9.I0.I12.Bit;
        real_rf_data[12][24] = dut.datapath.I24.I9.I0.I12.Bit;
        real_rf_data[12][25] = dut.datapath.I25.I9.I0.I12.Bit;
        real_rf_data[12][26] = dut.datapath.I26.I9.I0.I12.Bit;
        real_rf_data[12][27] = dut.datapath.I27.I9.I0.I12.Bit;
        real_rf_data[12][28] = dut.datapath.I28.I9.I0.I12.Bit;
        real_rf_data[12][29] = dut.datapath.I29.I9.I0.I12.Bit;
        real_rf_data[12][30] = dut.datapath.I30.I9.I0.I12.Bit;
        real_rf_data[12][31] = dut.datapath.I31.I9.I0.I12.Bit;
        real_rf_data[13][0] = dut.datapath.I0.I9.I0.I13.Bit;
        real_rf_data[13][1] = dut.datapath.I1.I9.I0.I13.Bit;
        real_rf_data[13][2] = dut.datapath.I2.I9.I0.I13.Bit;
        real_rf_data[13][3] = dut.datapath.I3.I9.I0.I13.Bit;
        real_rf_data[13][4] = dut.datapath.I4.I9.I0.I13.Bit;
        real_rf_data[13][5] = dut.datapath.I5.I9.I0.I13.Bit;
        real_rf_data[13][6] = dut.datapath.I6.I9.I0.I13.Bit;
        real_rf_data[13][7] = dut.datapath.I7.I9.I0.I13.Bit;
        real_rf_data[13][8] = dut.datapath.I8.I9.I0.I13.Bit;
        real_rf_data[13][9] = dut.datapath.I9.I9.I0.I13.Bit;
        real_rf_data[13][10] = dut.datapath.I10.I9.I0.I13.Bit;
        real_rf_data[13][11] = dut.datapath.I11.I9.I0.I13.Bit;
        real_rf_data[13][12] = dut.datapath.I12.I9.I0.I13.Bit;
        real_rf_data[13][13] = dut.datapath.I13.I9.I0.I13.Bit;
        real_rf_data[13][14] = dut.datapath.I14.I9.I0.I13.Bit;
        real_rf_data[13][15] = dut.datapath.I15.I9.I0.I13.Bit;
        real_rf_data[13][16] = dut.datapath.I16.I9.I0.I13.Bit;
        real_rf_data[13][17] = dut.datapath.I17.I9.I0.I13.Bit;
        real_rf_data[13][18] = dut.datapath.I18.I9.I0.I13.Bit;
        real_rf_data[13][19] = dut.datapath.I19.I9.I0.I13.Bit;
        real_rf_data[13][20] = dut.datapath.I20.I9.I0.I13.Bit;
        real_rf_data[13][21] = dut.datapath.I21.I9.I0.I13.Bit;
        real_rf_data[13][22] = dut.datapath.I22.I9.I0.I13.Bit;
        real_rf_data[13][23] = dut.datapath.I23.I9.I0.I13.Bit;
        real_rf_data[13][24] = dut.datapath.I24.I9.I0.I13.Bit;
        real_rf_data[13][25] = dut.datapath.I25.I9.I0.I13.Bit;
        real_rf_data[13][26] = dut.datapath.I26.I9.I0.I13.Bit;
        real_rf_data[13][27] = dut.datapath.I27.I9.I0.I13.Bit;
        real_rf_data[13][28] = dut.datapath.I28.I9.I0.I13.Bit;
        real_rf_data[13][29] = dut.datapath.I29.I9.I0.I13.Bit;
        real_rf_data[13][30] = dut.datapath.I30.I9.I0.I13.Bit;
        real_rf_data[13][31] = dut.datapath.I31.I9.I0.I13.Bit;
        real_rf_data[14][0] = dut.datapath.I0.I9.I0.I14.Bit;
        real_rf_data[14][1] = dut.datapath.I1.I9.I0.I14.Bit;
        real_rf_data[14][2] = dut.datapath.I2.I9.I0.I14.Bit;
        real_rf_data[14][3] = dut.datapath.I3.I9.I0.I14.Bit;
        real_rf_data[14][4] = dut.datapath.I4.I9.I0.I14.Bit;
        real_rf_data[14][5] = dut.datapath.I5.I9.I0.I14.Bit;
        real_rf_data[14][6] = dut.datapath.I6.I9.I0.I14.Bit;
        real_rf_data[14][7] = dut.datapath.I7.I9.I0.I14.Bit;
        real_rf_data[14][8] = dut.datapath.I8.I9.I0.I14.Bit;
        real_rf_data[14][9] = dut.datapath.I9.I9.I0.I14.Bit;
        real_rf_data[14][10] = dut.datapath.I10.I9.I0.I14.Bit;
        real_rf_data[14][11] = dut.datapath.I11.I9.I0.I14.Bit;
        real_rf_data[14][12] = dut.datapath.I12.I9.I0.I14.Bit;
        real_rf_data[14][13] = dut.datapath.I13.I9.I0.I14.Bit;
        real_rf_data[14][14] = dut.datapath.I14.I9.I0.I14.Bit;
        real_rf_data[14][15] = dut.datapath.I15.I9.I0.I14.Bit;
        real_rf_data[14][16] = dut.datapath.I16.I9.I0.I14.Bit;
        real_rf_data[14][17] = dut.datapath.I17.I9.I0.I14.Bit;
        real_rf_data[14][18] = dut.datapath.I18.I9.I0.I14.Bit;
        real_rf_data[14][19] = dut.datapath.I19.I9.I0.I14.Bit;
        real_rf_data[14][20] = dut.datapath.I20.I9.I0.I14.Bit;
        real_rf_data[14][21] = dut.datapath.I21.I9.I0.I14.Bit;
        real_rf_data[14][22] = dut.datapath.I22.I9.I0.I14.Bit;
        real_rf_data[14][23] = dut.datapath.I23.I9.I0.I14.Bit;
        real_rf_data[14][24] = dut.datapath.I24.I9.I0.I14.Bit;
        real_rf_data[14][25] = dut.datapath.I25.I9.I0.I14.Bit;
        real_rf_data[14][26] = dut.datapath.I26.I9.I0.I14.Bit;
        real_rf_data[14][27] = dut.datapath.I27.I9.I0.I14.Bit;
        real_rf_data[14][28] = dut.datapath.I28.I9.I0.I14.Bit;
        real_rf_data[14][29] = dut.datapath.I29.I9.I0.I14.Bit;
        real_rf_data[14][30] = dut.datapath.I30.I9.I0.I14.Bit;
        real_rf_data[14][31] = dut.datapath.I31.I9.I0.I14.Bit;
        real_rf_data[15][0] = dut.datapath.I0.I9.I0.I15.Bit;
        real_rf_data[15][1] = dut.datapath.I1.I9.I0.I15.Bit;
        real_rf_data[15][2] = dut.datapath.I2.I9.I0.I15.Bit;
        real_rf_data[15][3] = dut.datapath.I3.I9.I0.I15.Bit;
        real_rf_data[15][4] = dut.datapath.I4.I9.I0.I15.Bit;
        real_rf_data[15][5] = dut.datapath.I5.I9.I0.I15.Bit;
        real_rf_data[15][6] = dut.datapath.I6.I9.I0.I15.Bit;
        real_rf_data[15][7] = dut.datapath.I7.I9.I0.I15.Bit;
        real_rf_data[15][8] = dut.datapath.I8.I9.I0.I15.Bit;
        real_rf_data[15][9] = dut.datapath.I9.I9.I0.I15.Bit;
        real_rf_data[15][10] = dut.datapath.I10.I9.I0.I15.Bit;
        real_rf_data[15][11] = dut.datapath.I11.I9.I0.I15.Bit;
        real_rf_data[15][12] = dut.datapath.I12.I9.I0.I15.Bit;
        real_rf_data[15][13] = dut.datapath.I13.I9.I0.I15.Bit;
        real_rf_data[15][14] = dut.datapath.I14.I9.I0.I15.Bit;
        real_rf_data[15][15] = dut.datapath.I15.I9.I0.I15.Bit;
        real_rf_data[15][16] = dut.datapath.I16.I9.I0.I15.Bit;
        real_rf_data[15][17] = dut.datapath.I17.I9.I0.I15.Bit;
        real_rf_data[15][18] = dut.datapath.I18.I9.I0.I15.Bit;
        real_rf_data[15][19] = dut.datapath.I19.I9.I0.I15.Bit;
        real_rf_data[15][20] = dut.datapath.I20.I9.I0.I15.Bit;
        real_rf_data[15][21] = dut.datapath.I21.I9.I0.I15.Bit;
        real_rf_data[15][22] = dut.datapath.I22.I9.I0.I15.Bit;
        real_rf_data[15][23] = dut.datapath.I23.I9.I0.I15.Bit;
        real_rf_data[15][24] = dut.datapath.I24.I9.I0.I15.Bit;
        real_rf_data[15][25] = dut.datapath.I25.I9.I0.I15.Bit;
        real_rf_data[15][26] = dut.datapath.I26.I9.I0.I15.Bit;
        real_rf_data[15][27] = dut.datapath.I27.I9.I0.I15.Bit;
        real_rf_data[15][28] = dut.datapath.I28.I9.I0.I15.Bit;
        real_rf_data[15][29] = dut.datapath.I29.I9.I0.I15.Bit;
        real_rf_data[15][30] = dut.datapath.I30.I9.I0.I15.Bit;
        real_rf_data[15][31] = dut.datapath.I31.I9.I0.I15.Bit;
        real_rf_data[16][0] = dut.datapath.I0.I9.I0.I16.Bit;
        real_rf_data[16][1] = dut.datapath.I1.I9.I0.I16.Bit;
        real_rf_data[16][2] = dut.datapath.I2.I9.I0.I16.Bit;
        real_rf_data[16][3] = dut.datapath.I3.I9.I0.I16.Bit;
        real_rf_data[16][4] = dut.datapath.I4.I9.I0.I16.Bit;
        real_rf_data[16][5] = dut.datapath.I5.I9.I0.I16.Bit;
        real_rf_data[16][6] = dut.datapath.I6.I9.I0.I16.Bit;
        real_rf_data[16][7] = dut.datapath.I7.I9.I0.I16.Bit;
        real_rf_data[16][8] = dut.datapath.I8.I9.I0.I16.Bit;
        real_rf_data[16][9] = dut.datapath.I9.I9.I0.I16.Bit;
        real_rf_data[16][10] = dut.datapath.I10.I9.I0.I16.Bit;
        real_rf_data[16][11] = dut.datapath.I11.I9.I0.I16.Bit;
        real_rf_data[16][12] = dut.datapath.I12.I9.I0.I16.Bit;
        real_rf_data[16][13] = dut.datapath.I13.I9.I0.I16.Bit;
        real_rf_data[16][14] = dut.datapath.I14.I9.I0.I16.Bit;
        real_rf_data[16][15] = dut.datapath.I15.I9.I0.I16.Bit;
        real_rf_data[16][16] = dut.datapath.I16.I9.I0.I16.Bit;
        real_rf_data[16][17] = dut.datapath.I17.I9.I0.I16.Bit;
        real_rf_data[16][18] = dut.datapath.I18.I9.I0.I16.Bit;
        real_rf_data[16][19] = dut.datapath.I19.I9.I0.I16.Bit;
        real_rf_data[16][20] = dut.datapath.I20.I9.I0.I16.Bit;
        real_rf_data[16][21] = dut.datapath.I21.I9.I0.I16.Bit;
        real_rf_data[16][22] = dut.datapath.I22.I9.I0.I16.Bit;
        real_rf_data[16][23] = dut.datapath.I23.I9.I0.I16.Bit;
        real_rf_data[16][24] = dut.datapath.I24.I9.I0.I16.Bit;
        real_rf_data[16][25] = dut.datapath.I25.I9.I0.I16.Bit;
        real_rf_data[16][26] = dut.datapath.I26.I9.I0.I16.Bit;
        real_rf_data[16][27] = dut.datapath.I27.I9.I0.I16.Bit;
        real_rf_data[16][28] = dut.datapath.I28.I9.I0.I16.Bit;
        real_rf_data[16][29] = dut.datapath.I29.I9.I0.I16.Bit;
        real_rf_data[16][30] = dut.datapath.I30.I9.I0.I16.Bit;
        real_rf_data[16][31] = dut.datapath.I31.I9.I0.I16.Bit;
        real_rf_data[17][0] = dut.datapath.I0.I9.I0.I17.Bit;
        real_rf_data[17][1] = dut.datapath.I1.I9.I0.I17.Bit;
        real_rf_data[17][2] = dut.datapath.I2.I9.I0.I17.Bit;
        real_rf_data[17][3] = dut.datapath.I3.I9.I0.I17.Bit;
        real_rf_data[17][4] = dut.datapath.I4.I9.I0.I17.Bit;
        real_rf_data[17][5] = dut.datapath.I5.I9.I0.I17.Bit;
        real_rf_data[17][6] = dut.datapath.I6.I9.I0.I17.Bit;
        real_rf_data[17][7] = dut.datapath.I7.I9.I0.I17.Bit;
        real_rf_data[17][8] = dut.datapath.I8.I9.I0.I17.Bit;
        real_rf_data[17][9] = dut.datapath.I9.I9.I0.I17.Bit;
        real_rf_data[17][10] = dut.datapath.I10.I9.I0.I17.Bit;
        real_rf_data[17][11] = dut.datapath.I11.I9.I0.I17.Bit;
        real_rf_data[17][12] = dut.datapath.I12.I9.I0.I17.Bit;
        real_rf_data[17][13] = dut.datapath.I13.I9.I0.I17.Bit;
        real_rf_data[17][14] = dut.datapath.I14.I9.I0.I17.Bit;
        real_rf_data[17][15] = dut.datapath.I15.I9.I0.I17.Bit;
        real_rf_data[17][16] = dut.datapath.I16.I9.I0.I17.Bit;
        real_rf_data[17][17] = dut.datapath.I17.I9.I0.I17.Bit;
        real_rf_data[17][18] = dut.datapath.I18.I9.I0.I17.Bit;
        real_rf_data[17][19] = dut.datapath.I19.I9.I0.I17.Bit;
        real_rf_data[17][20] = dut.datapath.I20.I9.I0.I17.Bit;
        real_rf_data[17][21] = dut.datapath.I21.I9.I0.I17.Bit;
        real_rf_data[17][22] = dut.datapath.I22.I9.I0.I17.Bit;
        real_rf_data[17][23] = dut.datapath.I23.I9.I0.I17.Bit;
        real_rf_data[17][24] = dut.datapath.I24.I9.I0.I17.Bit;
        real_rf_data[17][25] = dut.datapath.I25.I9.I0.I17.Bit;
        real_rf_data[17][26] = dut.datapath.I26.I9.I0.I17.Bit;
        real_rf_data[17][27] = dut.datapath.I27.I9.I0.I17.Bit;
        real_rf_data[17][28] = dut.datapath.I28.I9.I0.I17.Bit;
        real_rf_data[17][29] = dut.datapath.I29.I9.I0.I17.Bit;
        real_rf_data[17][30] = dut.datapath.I30.I9.I0.I17.Bit;
        real_rf_data[17][31] = dut.datapath.I31.I9.I0.I17.Bit;
        real_rf_data[18][0] = dut.datapath.I0.I9.I0.I18.Bit;
        real_rf_data[18][1] = dut.datapath.I1.I9.I0.I18.Bit;
        real_rf_data[18][2] = dut.datapath.I2.I9.I0.I18.Bit;
        real_rf_data[18][3] = dut.datapath.I3.I9.I0.I18.Bit;
        real_rf_data[18][4] = dut.datapath.I4.I9.I0.I18.Bit;
        real_rf_data[18][5] = dut.datapath.I5.I9.I0.I18.Bit;
        real_rf_data[18][6] = dut.datapath.I6.I9.I0.I18.Bit;
        real_rf_data[18][7] = dut.datapath.I7.I9.I0.I18.Bit;
        real_rf_data[18][8] = dut.datapath.I8.I9.I0.I18.Bit;
        real_rf_data[18][9] = dut.datapath.I9.I9.I0.I18.Bit;
        real_rf_data[18][10] = dut.datapath.I10.I9.I0.I18.Bit;
        real_rf_data[18][11] = dut.datapath.I11.I9.I0.I18.Bit;
        real_rf_data[18][12] = dut.datapath.I12.I9.I0.I18.Bit;
        real_rf_data[18][13] = dut.datapath.I13.I9.I0.I18.Bit;
        real_rf_data[18][14] = dut.datapath.I14.I9.I0.I18.Bit;
        real_rf_data[18][15] = dut.datapath.I15.I9.I0.I18.Bit;
        real_rf_data[18][16] = dut.datapath.I16.I9.I0.I18.Bit;
        real_rf_data[18][17] = dut.datapath.I17.I9.I0.I18.Bit;
        real_rf_data[18][18] = dut.datapath.I18.I9.I0.I18.Bit;
        real_rf_data[18][19] = dut.datapath.I19.I9.I0.I18.Bit;
        real_rf_data[18][20] = dut.datapath.I20.I9.I0.I18.Bit;
        real_rf_data[18][21] = dut.datapath.I21.I9.I0.I18.Bit;
        real_rf_data[18][22] = dut.datapath.I22.I9.I0.I18.Bit;
        real_rf_data[18][23] = dut.datapath.I23.I9.I0.I18.Bit;
        real_rf_data[18][24] = dut.datapath.I24.I9.I0.I18.Bit;
        real_rf_data[18][25] = dut.datapath.I25.I9.I0.I18.Bit;
        real_rf_data[18][26] = dut.datapath.I26.I9.I0.I18.Bit;
        real_rf_data[18][27] = dut.datapath.I27.I9.I0.I18.Bit;
        real_rf_data[18][28] = dut.datapath.I28.I9.I0.I18.Bit;
        real_rf_data[18][29] = dut.datapath.I29.I9.I0.I18.Bit;
        real_rf_data[18][30] = dut.datapath.I30.I9.I0.I18.Bit;
        real_rf_data[18][31] = dut.datapath.I31.I9.I0.I18.Bit;
        real_rf_data[19][0] = dut.datapath.I0.I9.I0.I19.Bit;
        real_rf_data[19][1] = dut.datapath.I1.I9.I0.I19.Bit;
        real_rf_data[19][2] = dut.datapath.I2.I9.I0.I19.Bit;
        real_rf_data[19][3] = dut.datapath.I3.I9.I0.I19.Bit;
        real_rf_data[19][4] = dut.datapath.I4.I9.I0.I19.Bit;
        real_rf_data[19][5] = dut.datapath.I5.I9.I0.I19.Bit;
        real_rf_data[19][6] = dut.datapath.I6.I9.I0.I19.Bit;
        real_rf_data[19][7] = dut.datapath.I7.I9.I0.I19.Bit;
        real_rf_data[19][8] = dut.datapath.I8.I9.I0.I19.Bit;
        real_rf_data[19][9] = dut.datapath.I9.I9.I0.I19.Bit;
        real_rf_data[19][10] = dut.datapath.I10.I9.I0.I19.Bit;
        real_rf_data[19][11] = dut.datapath.I11.I9.I0.I19.Bit;
        real_rf_data[19][12] = dut.datapath.I12.I9.I0.I19.Bit;
        real_rf_data[19][13] = dut.datapath.I13.I9.I0.I19.Bit;
        real_rf_data[19][14] = dut.datapath.I14.I9.I0.I19.Bit;
        real_rf_data[19][15] = dut.datapath.I15.I9.I0.I19.Bit;
        real_rf_data[19][16] = dut.datapath.I16.I9.I0.I19.Bit;
        real_rf_data[19][17] = dut.datapath.I17.I9.I0.I19.Bit;
        real_rf_data[19][18] = dut.datapath.I18.I9.I0.I19.Bit;
        real_rf_data[19][19] = dut.datapath.I19.I9.I0.I19.Bit;
        real_rf_data[19][20] = dut.datapath.I20.I9.I0.I19.Bit;
        real_rf_data[19][21] = dut.datapath.I21.I9.I0.I19.Bit;
        real_rf_data[19][22] = dut.datapath.I22.I9.I0.I19.Bit;
        real_rf_data[19][23] = dut.datapath.I23.I9.I0.I19.Bit;
        real_rf_data[19][24] = dut.datapath.I24.I9.I0.I19.Bit;
        real_rf_data[19][25] = dut.datapath.I25.I9.I0.I19.Bit;
        real_rf_data[19][26] = dut.datapath.I26.I9.I0.I19.Bit;
        real_rf_data[19][27] = dut.datapath.I27.I9.I0.I19.Bit;
        real_rf_data[19][28] = dut.datapath.I28.I9.I0.I19.Bit;
        real_rf_data[19][29] = dut.datapath.I29.I9.I0.I19.Bit;
        real_rf_data[19][30] = dut.datapath.I30.I9.I0.I19.Bit;
        real_rf_data[19][31] = dut.datapath.I31.I9.I0.I19.Bit;
        real_rf_data[20][0] = dut.datapath.I0.I9.I0.I20.Bit;
        real_rf_data[20][1] = dut.datapath.I1.I9.I0.I20.Bit;
        real_rf_data[20][2] = dut.datapath.I2.I9.I0.I20.Bit;
        real_rf_data[20][3] = dut.datapath.I3.I9.I0.I20.Bit;
        real_rf_data[20][4] = dut.datapath.I4.I9.I0.I20.Bit;
        real_rf_data[20][5] = dut.datapath.I5.I9.I0.I20.Bit;
        real_rf_data[20][6] = dut.datapath.I6.I9.I0.I20.Bit;
        real_rf_data[20][7] = dut.datapath.I7.I9.I0.I20.Bit;
        real_rf_data[20][8] = dut.datapath.I8.I9.I0.I20.Bit;
        real_rf_data[20][9] = dut.datapath.I9.I9.I0.I20.Bit;
        real_rf_data[20][10] = dut.datapath.I10.I9.I0.I20.Bit;
        real_rf_data[20][11] = dut.datapath.I11.I9.I0.I20.Bit;
        real_rf_data[20][12] = dut.datapath.I12.I9.I0.I20.Bit;
        real_rf_data[20][13] = dut.datapath.I13.I9.I0.I20.Bit;
        real_rf_data[20][14] = dut.datapath.I14.I9.I0.I20.Bit;
        real_rf_data[20][15] = dut.datapath.I15.I9.I0.I20.Bit;
        real_rf_data[20][16] = dut.datapath.I16.I9.I0.I20.Bit;
        real_rf_data[20][17] = dut.datapath.I17.I9.I0.I20.Bit;
        real_rf_data[20][18] = dut.datapath.I18.I9.I0.I20.Bit;
        real_rf_data[20][19] = dut.datapath.I19.I9.I0.I20.Bit;
        real_rf_data[20][20] = dut.datapath.I20.I9.I0.I20.Bit;
        real_rf_data[20][21] = dut.datapath.I21.I9.I0.I20.Bit;
        real_rf_data[20][22] = dut.datapath.I22.I9.I0.I20.Bit;
        real_rf_data[20][23] = dut.datapath.I23.I9.I0.I20.Bit;
        real_rf_data[20][24] = dut.datapath.I24.I9.I0.I20.Bit;
        real_rf_data[20][25] = dut.datapath.I25.I9.I0.I20.Bit;
        real_rf_data[20][26] = dut.datapath.I26.I9.I0.I20.Bit;
        real_rf_data[20][27] = dut.datapath.I27.I9.I0.I20.Bit;
        real_rf_data[20][28] = dut.datapath.I28.I9.I0.I20.Bit;
        real_rf_data[20][29] = dut.datapath.I29.I9.I0.I20.Bit;
        real_rf_data[20][30] = dut.datapath.I30.I9.I0.I20.Bit;
        real_rf_data[20][31] = dut.datapath.I31.I9.I0.I20.Bit;
        real_rf_data[21][0] = dut.datapath.I0.I9.I0.I21.Bit;
        real_rf_data[21][1] = dut.datapath.I1.I9.I0.I21.Bit;
        real_rf_data[21][2] = dut.datapath.I2.I9.I0.I21.Bit;
        real_rf_data[21][3] = dut.datapath.I3.I9.I0.I21.Bit;
        real_rf_data[21][4] = dut.datapath.I4.I9.I0.I21.Bit;
        real_rf_data[21][5] = dut.datapath.I5.I9.I0.I21.Bit;
        real_rf_data[21][6] = dut.datapath.I6.I9.I0.I21.Bit;
        real_rf_data[21][7] = dut.datapath.I7.I9.I0.I21.Bit;
        real_rf_data[21][8] = dut.datapath.I8.I9.I0.I21.Bit;
        real_rf_data[21][9] = dut.datapath.I9.I9.I0.I21.Bit;
        real_rf_data[21][10] = dut.datapath.I10.I9.I0.I21.Bit;
        real_rf_data[21][11] = dut.datapath.I11.I9.I0.I21.Bit;
        real_rf_data[21][12] = dut.datapath.I12.I9.I0.I21.Bit;
        real_rf_data[21][13] = dut.datapath.I13.I9.I0.I21.Bit;
        real_rf_data[21][14] = dut.datapath.I14.I9.I0.I21.Bit;
        real_rf_data[21][15] = dut.datapath.I15.I9.I0.I21.Bit;
        real_rf_data[21][16] = dut.datapath.I16.I9.I0.I21.Bit;
        real_rf_data[21][17] = dut.datapath.I17.I9.I0.I21.Bit;
        real_rf_data[21][18] = dut.datapath.I18.I9.I0.I21.Bit;
        real_rf_data[21][19] = dut.datapath.I19.I9.I0.I21.Bit;
        real_rf_data[21][20] = dut.datapath.I20.I9.I0.I21.Bit;
        real_rf_data[21][21] = dut.datapath.I21.I9.I0.I21.Bit;
        real_rf_data[21][22] = dut.datapath.I22.I9.I0.I21.Bit;
        real_rf_data[21][23] = dut.datapath.I23.I9.I0.I21.Bit;
        real_rf_data[21][24] = dut.datapath.I24.I9.I0.I21.Bit;
        real_rf_data[21][25] = dut.datapath.I25.I9.I0.I21.Bit;
        real_rf_data[21][26] = dut.datapath.I26.I9.I0.I21.Bit;
        real_rf_data[21][27] = dut.datapath.I27.I9.I0.I21.Bit;
        real_rf_data[21][28] = dut.datapath.I28.I9.I0.I21.Bit;
        real_rf_data[21][29] = dut.datapath.I29.I9.I0.I21.Bit;
        real_rf_data[21][30] = dut.datapath.I30.I9.I0.I21.Bit;
        real_rf_data[21][31] = dut.datapath.I31.I9.I0.I21.Bit;
        real_rf_data[22][0] = dut.datapath.I0.I9.I0.I22.Bit;
        real_rf_data[22][1] = dut.datapath.I1.I9.I0.I22.Bit;
        real_rf_data[22][2] = dut.datapath.I2.I9.I0.I22.Bit;
        real_rf_data[22][3] = dut.datapath.I3.I9.I0.I22.Bit;
        real_rf_data[22][4] = dut.datapath.I4.I9.I0.I22.Bit;
        real_rf_data[22][5] = dut.datapath.I5.I9.I0.I22.Bit;
        real_rf_data[22][6] = dut.datapath.I6.I9.I0.I22.Bit;
        real_rf_data[22][7] = dut.datapath.I7.I9.I0.I22.Bit;
        real_rf_data[22][8] = dut.datapath.I8.I9.I0.I22.Bit;
        real_rf_data[22][9] = dut.datapath.I9.I9.I0.I22.Bit;
        real_rf_data[22][10] = dut.datapath.I10.I9.I0.I22.Bit;
        real_rf_data[22][11] = dut.datapath.I11.I9.I0.I22.Bit;
        real_rf_data[22][12] = dut.datapath.I12.I9.I0.I22.Bit;
        real_rf_data[22][13] = dut.datapath.I13.I9.I0.I22.Bit;
        real_rf_data[22][14] = dut.datapath.I14.I9.I0.I22.Bit;
        real_rf_data[22][15] = dut.datapath.I15.I9.I0.I22.Bit;
        real_rf_data[22][16] = dut.datapath.I16.I9.I0.I22.Bit;
        real_rf_data[22][17] = dut.datapath.I17.I9.I0.I22.Bit;
        real_rf_data[22][18] = dut.datapath.I18.I9.I0.I22.Bit;
        real_rf_data[22][19] = dut.datapath.I19.I9.I0.I22.Bit;
        real_rf_data[22][20] = dut.datapath.I20.I9.I0.I22.Bit;
        real_rf_data[22][21] = dut.datapath.I21.I9.I0.I22.Bit;
        real_rf_data[22][22] = dut.datapath.I22.I9.I0.I22.Bit;
        real_rf_data[22][23] = dut.datapath.I23.I9.I0.I22.Bit;
        real_rf_data[22][24] = dut.datapath.I24.I9.I0.I22.Bit;
        real_rf_data[22][25] = dut.datapath.I25.I9.I0.I22.Bit;
        real_rf_data[22][26] = dut.datapath.I26.I9.I0.I22.Bit;
        real_rf_data[22][27] = dut.datapath.I27.I9.I0.I22.Bit;
        real_rf_data[22][28] = dut.datapath.I28.I9.I0.I22.Bit;
        real_rf_data[22][29] = dut.datapath.I29.I9.I0.I22.Bit;
        real_rf_data[22][30] = dut.datapath.I30.I9.I0.I22.Bit;
        real_rf_data[22][31] = dut.datapath.I31.I9.I0.I22.Bit;
        real_rf_data[23][0] = dut.datapath.I0.I9.I0.I23.Bit;
        real_rf_data[23][1] = dut.datapath.I1.I9.I0.I23.Bit;
        real_rf_data[23][2] = dut.datapath.I2.I9.I0.I23.Bit;
        real_rf_data[23][3] = dut.datapath.I3.I9.I0.I23.Bit;
        real_rf_data[23][4] = dut.datapath.I4.I9.I0.I23.Bit;
        real_rf_data[23][5] = dut.datapath.I5.I9.I0.I23.Bit;
        real_rf_data[23][6] = dut.datapath.I6.I9.I0.I23.Bit;
        real_rf_data[23][7] = dut.datapath.I7.I9.I0.I23.Bit;
        real_rf_data[23][8] = dut.datapath.I8.I9.I0.I23.Bit;
        real_rf_data[23][9] = dut.datapath.I9.I9.I0.I23.Bit;
        real_rf_data[23][10] = dut.datapath.I10.I9.I0.I23.Bit;
        real_rf_data[23][11] = dut.datapath.I11.I9.I0.I23.Bit;
        real_rf_data[23][12] = dut.datapath.I12.I9.I0.I23.Bit;
        real_rf_data[23][13] = dut.datapath.I13.I9.I0.I23.Bit;
        real_rf_data[23][14] = dut.datapath.I14.I9.I0.I23.Bit;
        real_rf_data[23][15] = dut.datapath.I15.I9.I0.I23.Bit;
        real_rf_data[23][16] = dut.datapath.I16.I9.I0.I23.Bit;
        real_rf_data[23][17] = dut.datapath.I17.I9.I0.I23.Bit;
        real_rf_data[23][18] = dut.datapath.I18.I9.I0.I23.Bit;
        real_rf_data[23][19] = dut.datapath.I19.I9.I0.I23.Bit;
        real_rf_data[23][20] = dut.datapath.I20.I9.I0.I23.Bit;
        real_rf_data[23][21] = dut.datapath.I21.I9.I0.I23.Bit;
        real_rf_data[23][22] = dut.datapath.I22.I9.I0.I23.Bit;
        real_rf_data[23][23] = dut.datapath.I23.I9.I0.I23.Bit;
        real_rf_data[23][24] = dut.datapath.I24.I9.I0.I23.Bit;
        real_rf_data[23][25] = dut.datapath.I25.I9.I0.I23.Bit;
        real_rf_data[23][26] = dut.datapath.I26.I9.I0.I23.Bit;
        real_rf_data[23][27] = dut.datapath.I27.I9.I0.I23.Bit;
        real_rf_data[23][28] = dut.datapath.I28.I9.I0.I23.Bit;
        real_rf_data[23][29] = dut.datapath.I29.I9.I0.I23.Bit;
        real_rf_data[23][30] = dut.datapath.I30.I9.I0.I23.Bit;
        real_rf_data[23][31] = dut.datapath.I31.I9.I0.I23.Bit;
        real_rf_data[24][0] = dut.datapath.I0.I9.I0.I24.Bit;
        real_rf_data[24][1] = dut.datapath.I1.I9.I0.I24.Bit;
        real_rf_data[24][2] = dut.datapath.I2.I9.I0.I24.Bit;
        real_rf_data[24][3] = dut.datapath.I3.I9.I0.I24.Bit;
        real_rf_data[24][4] = dut.datapath.I4.I9.I0.I24.Bit;
        real_rf_data[24][5] = dut.datapath.I5.I9.I0.I24.Bit;
        real_rf_data[24][6] = dut.datapath.I6.I9.I0.I24.Bit;
        real_rf_data[24][7] = dut.datapath.I7.I9.I0.I24.Bit;
        real_rf_data[24][8] = dut.datapath.I8.I9.I0.I24.Bit;
        real_rf_data[24][9] = dut.datapath.I9.I9.I0.I24.Bit;
        real_rf_data[24][10] = dut.datapath.I10.I9.I0.I24.Bit;
        real_rf_data[24][11] = dut.datapath.I11.I9.I0.I24.Bit;
        real_rf_data[24][12] = dut.datapath.I12.I9.I0.I24.Bit;
        real_rf_data[24][13] = dut.datapath.I13.I9.I0.I24.Bit;
        real_rf_data[24][14] = dut.datapath.I14.I9.I0.I24.Bit;
        real_rf_data[24][15] = dut.datapath.I15.I9.I0.I24.Bit;
        real_rf_data[24][16] = dut.datapath.I16.I9.I0.I24.Bit;
        real_rf_data[24][17] = dut.datapath.I17.I9.I0.I24.Bit;
        real_rf_data[24][18] = dut.datapath.I18.I9.I0.I24.Bit;
        real_rf_data[24][19] = dut.datapath.I19.I9.I0.I24.Bit;
        real_rf_data[24][20] = dut.datapath.I20.I9.I0.I24.Bit;
        real_rf_data[24][21] = dut.datapath.I21.I9.I0.I24.Bit;
        real_rf_data[24][22] = dut.datapath.I22.I9.I0.I24.Bit;
        real_rf_data[24][23] = dut.datapath.I23.I9.I0.I24.Bit;
        real_rf_data[24][24] = dut.datapath.I24.I9.I0.I24.Bit;
        real_rf_data[24][25] = dut.datapath.I25.I9.I0.I24.Bit;
        real_rf_data[24][26] = dut.datapath.I26.I9.I0.I24.Bit;
        real_rf_data[24][27] = dut.datapath.I27.I9.I0.I24.Bit;
        real_rf_data[24][28] = dut.datapath.I28.I9.I0.I24.Bit;
        real_rf_data[24][29] = dut.datapath.I29.I9.I0.I24.Bit;
        real_rf_data[24][30] = dut.datapath.I30.I9.I0.I24.Bit;
        real_rf_data[24][31] = dut.datapath.I31.I9.I0.I24.Bit;
        real_rf_data[25][0] = dut.datapath.I0.I9.I0.I25.Bit;
        real_rf_data[25][1] = dut.datapath.I1.I9.I0.I25.Bit;
        real_rf_data[25][2] = dut.datapath.I2.I9.I0.I25.Bit;
        real_rf_data[25][3] = dut.datapath.I3.I9.I0.I25.Bit;
        real_rf_data[25][4] = dut.datapath.I4.I9.I0.I25.Bit;
        real_rf_data[25][5] = dut.datapath.I5.I9.I0.I25.Bit;
        real_rf_data[25][6] = dut.datapath.I6.I9.I0.I25.Bit;
        real_rf_data[25][7] = dut.datapath.I7.I9.I0.I25.Bit;
        real_rf_data[25][8] = dut.datapath.I8.I9.I0.I25.Bit;
        real_rf_data[25][9] = dut.datapath.I9.I9.I0.I25.Bit;
        real_rf_data[25][10] = dut.datapath.I10.I9.I0.I25.Bit;
        real_rf_data[25][11] = dut.datapath.I11.I9.I0.I25.Bit;
        real_rf_data[25][12] = dut.datapath.I12.I9.I0.I25.Bit;
        real_rf_data[25][13] = dut.datapath.I13.I9.I0.I25.Bit;
        real_rf_data[25][14] = dut.datapath.I14.I9.I0.I25.Bit;
        real_rf_data[25][15] = dut.datapath.I15.I9.I0.I25.Bit;
        real_rf_data[25][16] = dut.datapath.I16.I9.I0.I25.Bit;
        real_rf_data[25][17] = dut.datapath.I17.I9.I0.I25.Bit;
        real_rf_data[25][18] = dut.datapath.I18.I9.I0.I25.Bit;
        real_rf_data[25][19] = dut.datapath.I19.I9.I0.I25.Bit;
        real_rf_data[25][20] = dut.datapath.I20.I9.I0.I25.Bit;
        real_rf_data[25][21] = dut.datapath.I21.I9.I0.I25.Bit;
        real_rf_data[25][22] = dut.datapath.I22.I9.I0.I25.Bit;
        real_rf_data[25][23] = dut.datapath.I23.I9.I0.I25.Bit;
        real_rf_data[25][24] = dut.datapath.I24.I9.I0.I25.Bit;
        real_rf_data[25][25] = dut.datapath.I25.I9.I0.I25.Bit;
        real_rf_data[25][26] = dut.datapath.I26.I9.I0.I25.Bit;
        real_rf_data[25][27] = dut.datapath.I27.I9.I0.I25.Bit;
        real_rf_data[25][28] = dut.datapath.I28.I9.I0.I25.Bit;
        real_rf_data[25][29] = dut.datapath.I29.I9.I0.I25.Bit;
        real_rf_data[25][30] = dut.datapath.I30.I9.I0.I25.Bit;
        real_rf_data[25][31] = dut.datapath.I31.I9.I0.I25.Bit;
        real_rf_data[26][0] = dut.datapath.I0.I9.I0.I26.Bit;
        real_rf_data[26][1] = dut.datapath.I1.I9.I0.I26.Bit;
        real_rf_data[26][2] = dut.datapath.I2.I9.I0.I26.Bit;
        real_rf_data[26][3] = dut.datapath.I3.I9.I0.I26.Bit;
        real_rf_data[26][4] = dut.datapath.I4.I9.I0.I26.Bit;
        real_rf_data[26][5] = dut.datapath.I5.I9.I0.I26.Bit;
        real_rf_data[26][6] = dut.datapath.I6.I9.I0.I26.Bit;
        real_rf_data[26][7] = dut.datapath.I7.I9.I0.I26.Bit;
        real_rf_data[26][8] = dut.datapath.I8.I9.I0.I26.Bit;
        real_rf_data[26][9] = dut.datapath.I9.I9.I0.I26.Bit;
        real_rf_data[26][10] = dut.datapath.I10.I9.I0.I26.Bit;
        real_rf_data[26][11] = dut.datapath.I11.I9.I0.I26.Bit;
        real_rf_data[26][12] = dut.datapath.I12.I9.I0.I26.Bit;
        real_rf_data[26][13] = dut.datapath.I13.I9.I0.I26.Bit;
        real_rf_data[26][14] = dut.datapath.I14.I9.I0.I26.Bit;
        real_rf_data[26][15] = dut.datapath.I15.I9.I0.I26.Bit;
        real_rf_data[26][16] = dut.datapath.I16.I9.I0.I26.Bit;
        real_rf_data[26][17] = dut.datapath.I17.I9.I0.I26.Bit;
        real_rf_data[26][18] = dut.datapath.I18.I9.I0.I26.Bit;
        real_rf_data[26][19] = dut.datapath.I19.I9.I0.I26.Bit;
        real_rf_data[26][20] = dut.datapath.I20.I9.I0.I26.Bit;
        real_rf_data[26][21] = dut.datapath.I21.I9.I0.I26.Bit;
        real_rf_data[26][22] = dut.datapath.I22.I9.I0.I26.Bit;
        real_rf_data[26][23] = dut.datapath.I23.I9.I0.I26.Bit;
        real_rf_data[26][24] = dut.datapath.I24.I9.I0.I26.Bit;
        real_rf_data[26][25] = dut.datapath.I25.I9.I0.I26.Bit;
        real_rf_data[26][26] = dut.datapath.I26.I9.I0.I26.Bit;
        real_rf_data[26][27] = dut.datapath.I27.I9.I0.I26.Bit;
        real_rf_data[26][28] = dut.datapath.I28.I9.I0.I26.Bit;
        real_rf_data[26][29] = dut.datapath.I29.I9.I0.I26.Bit;
        real_rf_data[26][30] = dut.datapath.I30.I9.I0.I26.Bit;
        real_rf_data[26][31] = dut.datapath.I31.I9.I0.I26.Bit;
        real_rf_data[27][0] = dut.datapath.I0.I9.I0.I27.Bit;
        real_rf_data[27][1] = dut.datapath.I1.I9.I0.I27.Bit;
        real_rf_data[27][2] = dut.datapath.I2.I9.I0.I27.Bit;
        real_rf_data[27][3] = dut.datapath.I3.I9.I0.I27.Bit;
        real_rf_data[27][4] = dut.datapath.I4.I9.I0.I27.Bit;
        real_rf_data[27][5] = dut.datapath.I5.I9.I0.I27.Bit;
        real_rf_data[27][6] = dut.datapath.I6.I9.I0.I27.Bit;
        real_rf_data[27][7] = dut.datapath.I7.I9.I0.I27.Bit;
        real_rf_data[27][8] = dut.datapath.I8.I9.I0.I27.Bit;
        real_rf_data[27][9] = dut.datapath.I9.I9.I0.I27.Bit;
        real_rf_data[27][10] = dut.datapath.I10.I9.I0.I27.Bit;
        real_rf_data[27][11] = dut.datapath.I11.I9.I0.I27.Bit;
        real_rf_data[27][12] = dut.datapath.I12.I9.I0.I27.Bit;
        real_rf_data[27][13] = dut.datapath.I13.I9.I0.I27.Bit;
        real_rf_data[27][14] = dut.datapath.I14.I9.I0.I27.Bit;
        real_rf_data[27][15] = dut.datapath.I15.I9.I0.I27.Bit;
        real_rf_data[27][16] = dut.datapath.I16.I9.I0.I27.Bit;
        real_rf_data[27][17] = dut.datapath.I17.I9.I0.I27.Bit;
        real_rf_data[27][18] = dut.datapath.I18.I9.I0.I27.Bit;
        real_rf_data[27][19] = dut.datapath.I19.I9.I0.I27.Bit;
        real_rf_data[27][20] = dut.datapath.I20.I9.I0.I27.Bit;
        real_rf_data[27][21] = dut.datapath.I21.I9.I0.I27.Bit;
        real_rf_data[27][22] = dut.datapath.I22.I9.I0.I27.Bit;
        real_rf_data[27][23] = dut.datapath.I23.I9.I0.I27.Bit;
        real_rf_data[27][24] = dut.datapath.I24.I9.I0.I27.Bit;
        real_rf_data[27][25] = dut.datapath.I25.I9.I0.I27.Bit;
        real_rf_data[27][26] = dut.datapath.I26.I9.I0.I27.Bit;
        real_rf_data[27][27] = dut.datapath.I27.I9.I0.I27.Bit;
        real_rf_data[27][28] = dut.datapath.I28.I9.I0.I27.Bit;
        real_rf_data[27][29] = dut.datapath.I29.I9.I0.I27.Bit;
        real_rf_data[27][30] = dut.datapath.I30.I9.I0.I27.Bit;
        real_rf_data[27][31] = dut.datapath.I31.I9.I0.I27.Bit;
        real_rf_data[28][0] = dut.datapath.I0.I9.I0.I28.Bit;
        real_rf_data[28][1] = dut.datapath.I1.I9.I0.I28.Bit;
        real_rf_data[28][2] = dut.datapath.I2.I9.I0.I28.Bit;
        real_rf_data[28][3] = dut.datapath.I3.I9.I0.I28.Bit;
        real_rf_data[28][4] = dut.datapath.I4.I9.I0.I28.Bit;
        real_rf_data[28][5] = dut.datapath.I5.I9.I0.I28.Bit;
        real_rf_data[28][6] = dut.datapath.I6.I9.I0.I28.Bit;
        real_rf_data[28][7] = dut.datapath.I7.I9.I0.I28.Bit;
        real_rf_data[28][8] = dut.datapath.I8.I9.I0.I28.Bit;
        real_rf_data[28][9] = dut.datapath.I9.I9.I0.I28.Bit;
        real_rf_data[28][10] = dut.datapath.I10.I9.I0.I28.Bit;
        real_rf_data[28][11] = dut.datapath.I11.I9.I0.I28.Bit;
        real_rf_data[28][12] = dut.datapath.I12.I9.I0.I28.Bit;
        real_rf_data[28][13] = dut.datapath.I13.I9.I0.I28.Bit;
        real_rf_data[28][14] = dut.datapath.I14.I9.I0.I28.Bit;
        real_rf_data[28][15] = dut.datapath.I15.I9.I0.I28.Bit;
        real_rf_data[28][16] = dut.datapath.I16.I9.I0.I28.Bit;
        real_rf_data[28][17] = dut.datapath.I17.I9.I0.I28.Bit;
        real_rf_data[28][18] = dut.datapath.I18.I9.I0.I28.Bit;
        real_rf_data[28][19] = dut.datapath.I19.I9.I0.I28.Bit;
        real_rf_data[28][20] = dut.datapath.I20.I9.I0.I28.Bit;
        real_rf_data[28][21] = dut.datapath.I21.I9.I0.I28.Bit;
        real_rf_data[28][22] = dut.datapath.I22.I9.I0.I28.Bit;
        real_rf_data[28][23] = dut.datapath.I23.I9.I0.I28.Bit;
        real_rf_data[28][24] = dut.datapath.I24.I9.I0.I28.Bit;
        real_rf_data[28][25] = dut.datapath.I25.I9.I0.I28.Bit;
        real_rf_data[28][26] = dut.datapath.I26.I9.I0.I28.Bit;
        real_rf_data[28][27] = dut.datapath.I27.I9.I0.I28.Bit;
        real_rf_data[28][28] = dut.datapath.I28.I9.I0.I28.Bit;
        real_rf_data[28][29] = dut.datapath.I29.I9.I0.I28.Bit;
        real_rf_data[28][30] = dut.datapath.I30.I9.I0.I28.Bit;
        real_rf_data[28][31] = dut.datapath.I31.I9.I0.I28.Bit;
        real_rf_data[29][0] = dut.datapath.I0.I9.I0.I29.Bit;
        real_rf_data[29][1] = dut.datapath.I1.I9.I0.I29.Bit;
        real_rf_data[29][2] = dut.datapath.I2.I9.I0.I29.Bit;
        real_rf_data[29][3] = dut.datapath.I3.I9.I0.I29.Bit;
        real_rf_data[29][4] = dut.datapath.I4.I9.I0.I29.Bit;
        real_rf_data[29][5] = dut.datapath.I5.I9.I0.I29.Bit;
        real_rf_data[29][6] = dut.datapath.I6.I9.I0.I29.Bit;
        real_rf_data[29][7] = dut.datapath.I7.I9.I0.I29.Bit;
        real_rf_data[29][8] = dut.datapath.I8.I9.I0.I29.Bit;
        real_rf_data[29][9] = dut.datapath.I9.I9.I0.I29.Bit;
        real_rf_data[29][10] = dut.datapath.I10.I9.I0.I29.Bit;
        real_rf_data[29][11] = dut.datapath.I11.I9.I0.I29.Bit;
        real_rf_data[29][12] = dut.datapath.I12.I9.I0.I29.Bit;
        real_rf_data[29][13] = dut.datapath.I13.I9.I0.I29.Bit;
        real_rf_data[29][14] = dut.datapath.I14.I9.I0.I29.Bit;
        real_rf_data[29][15] = dut.datapath.I15.I9.I0.I29.Bit;
        real_rf_data[29][16] = dut.datapath.I16.I9.I0.I29.Bit;
        real_rf_data[29][17] = dut.datapath.I17.I9.I0.I29.Bit;
        real_rf_data[29][18] = dut.datapath.I18.I9.I0.I29.Bit;
        real_rf_data[29][19] = dut.datapath.I19.I9.I0.I29.Bit;
        real_rf_data[29][20] = dut.datapath.I20.I9.I0.I29.Bit;
        real_rf_data[29][21] = dut.datapath.I21.I9.I0.I29.Bit;
        real_rf_data[29][22] = dut.datapath.I22.I9.I0.I29.Bit;
        real_rf_data[29][23] = dut.datapath.I23.I9.I0.I29.Bit;
        real_rf_data[29][24] = dut.datapath.I24.I9.I0.I29.Bit;
        real_rf_data[29][25] = dut.datapath.I25.I9.I0.I29.Bit;
        real_rf_data[29][26] = dut.datapath.I26.I9.I0.I29.Bit;
        real_rf_data[29][27] = dut.datapath.I27.I9.I0.I29.Bit;
        real_rf_data[29][28] = dut.datapath.I28.I9.I0.I29.Bit;
        real_rf_data[29][29] = dut.datapath.I29.I9.I0.I29.Bit;
        real_rf_data[29][30] = dut.datapath.I30.I9.I0.I29.Bit;
        real_rf_data[29][31] = dut.datapath.I31.I9.I0.I29.Bit;
        real_rf_data[30][0] = dut.datapath.I0.I9.I0.I30.Bit;
        real_rf_data[30][1] = dut.datapath.I1.I9.I0.I30.Bit;
        real_rf_data[30][2] = dut.datapath.I2.I9.I0.I30.Bit;
        real_rf_data[30][3] = dut.datapath.I3.I9.I0.I30.Bit;
        real_rf_data[30][4] = dut.datapath.I4.I9.I0.I30.Bit;
        real_rf_data[30][5] = dut.datapath.I5.I9.I0.I30.Bit;
        real_rf_data[30][6] = dut.datapath.I6.I9.I0.I30.Bit;
        real_rf_data[30][7] = dut.datapath.I7.I9.I0.I30.Bit;
        real_rf_data[30][8] = dut.datapath.I8.I9.I0.I30.Bit;
        real_rf_data[30][9] = dut.datapath.I9.I9.I0.I30.Bit;
        real_rf_data[30][10] = dut.datapath.I10.I9.I0.I30.Bit;
        real_rf_data[30][11] = dut.datapath.I11.I9.I0.I30.Bit;
        real_rf_data[30][12] = dut.datapath.I12.I9.I0.I30.Bit;
        real_rf_data[30][13] = dut.datapath.I13.I9.I0.I30.Bit;
        real_rf_data[30][14] = dut.datapath.I14.I9.I0.I30.Bit;
        real_rf_data[30][15] = dut.datapath.I15.I9.I0.I30.Bit;
        real_rf_data[30][16] = dut.datapath.I16.I9.I0.I30.Bit;
        real_rf_data[30][17] = dut.datapath.I17.I9.I0.I30.Bit;
        real_rf_data[30][18] = dut.datapath.I18.I9.I0.I30.Bit;
        real_rf_data[30][19] = dut.datapath.I19.I9.I0.I30.Bit;
        real_rf_data[30][20] = dut.datapath.I20.I9.I0.I30.Bit;
        real_rf_data[30][21] = dut.datapath.I21.I9.I0.I30.Bit;
        real_rf_data[30][22] = dut.datapath.I22.I9.I0.I30.Bit;
        real_rf_data[30][23] = dut.datapath.I23.I9.I0.I30.Bit;
        real_rf_data[30][24] = dut.datapath.I24.I9.I0.I30.Bit;
        real_rf_data[30][25] = dut.datapath.I25.I9.I0.I30.Bit;
        real_rf_data[30][26] = dut.datapath.I26.I9.I0.I30.Bit;
        real_rf_data[30][27] = dut.datapath.I27.I9.I0.I30.Bit;
        real_rf_data[30][28] = dut.datapath.I28.I9.I0.I30.Bit;
        real_rf_data[30][29] = dut.datapath.I29.I9.I0.I30.Bit;
        real_rf_data[30][30] = dut.datapath.I30.I9.I0.I30.Bit;
        real_rf_data[30][31] = dut.datapath.I31.I9.I0.I30.Bit;
        real_rf_data[31][0] = dut.datapath.I0.I9.I0.I31.Bit;
        real_rf_data[31][1] = dut.datapath.I1.I9.I0.I31.Bit;
        real_rf_data[31][2] = dut.datapath.I2.I9.I0.I31.Bit;
        real_rf_data[31][3] = dut.datapath.I3.I9.I0.I31.Bit;
        real_rf_data[31][4] = dut.datapath.I4.I9.I0.I31.Bit;
        real_rf_data[31][5] = dut.datapath.I5.I9.I0.I31.Bit;
        real_rf_data[31][6] = dut.datapath.I6.I9.I0.I31.Bit;
        real_rf_data[31][7] = dut.datapath.I7.I9.I0.I31.Bit;
        real_rf_data[31][8] = dut.datapath.I8.I9.I0.I31.Bit;
        real_rf_data[31][9] = dut.datapath.I9.I9.I0.I31.Bit;
        real_rf_data[31][10] = dut.datapath.I10.I9.I0.I31.Bit;
        real_rf_data[31][11] = dut.datapath.I11.I9.I0.I31.Bit;
        real_rf_data[31][12] = dut.datapath.I12.I9.I0.I31.Bit;
        real_rf_data[31][13] = dut.datapath.I13.I9.I0.I31.Bit;
        real_rf_data[31][14] = dut.datapath.I14.I9.I0.I31.Bit;
        real_rf_data[31][15] = dut.datapath.I15.I9.I0.I31.Bit;
        real_rf_data[31][16] = dut.datapath.I16.I9.I0.I31.Bit;
        real_rf_data[31][17] = dut.datapath.I17.I9.I0.I31.Bit;
        real_rf_data[31][18] = dut.datapath.I18.I9.I0.I31.Bit;
        real_rf_data[31][19] = dut.datapath.I19.I9.I0.I31.Bit;
        real_rf_data[31][20] = dut.datapath.I20.I9.I0.I31.Bit;
        real_rf_data[31][21] = dut.datapath.I21.I9.I0.I31.Bit;
        real_rf_data[31][22] = dut.datapath.I22.I9.I0.I31.Bit;
        real_rf_data[31][23] = dut.datapath.I23.I9.I0.I31.Bit;
        real_rf_data[31][24] = dut.datapath.I24.I9.I0.I31.Bit;
        real_rf_data[31][25] = dut.datapath.I25.I9.I0.I31.Bit;
        real_rf_data[31][26] = dut.datapath.I26.I9.I0.I31.Bit;
        real_rf_data[31][27] = dut.datapath.I27.I9.I0.I31.Bit;
        real_rf_data[31][28] = dut.datapath.I28.I9.I0.I31.Bit;
        real_rf_data[31][29] = dut.datapath.I29.I9.I0.I31.Bit;
        real_rf_data[31][30] = dut.datapath.I30.I9.I0.I31.Bit;
        real_rf_data[31][31] = dut.datapath.I31.I9.I0.I31.Bit;
    end

    always_comb begin
        mon_itf.valid       = ~rst;
        mon_itf.order       = '0;
        mon_itf.inst        = imem_rdata;
        mon_itf.rs1_addr    = dut.control.rs1_s;
        mon_itf.rs2_addr    = dut.control.rs2_s;
        mon_itf.rs1_rdata   = rs1_rdata;
        mon_itf.rs2_rdata   = dmem_wdata;
        mon_itf.rd_addr     = dut.control.rd_s;
        mon_itf.rd_wdata    = rd_wdata;
        mon_itf.pc_rdata    = imem_addr;
        mon_itf.pc_wdata    = pc_wdata;
        mon_itf.mem_addr    = dmem_addr;
        mon_itf.mem_rmask   = dut.control.dmem_rmask;
        mon_itf.mem_wmask   = dmem_wmask;
        mon_itf.mem_rdata   = dmem_rdata;
        mon_itf.mem_wdata   = dmem_wdata;
    end

    initial begin
        $fsdbDumpfile("dump.fsdb");
        $fsdbDumpvars(0, "+all");
        rst = 1'b1;
        repeat (2) @(posedge clk);
        rst <= 1'b0;
        #100000000;
        $finish;
    end

endmodule
