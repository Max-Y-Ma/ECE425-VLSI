* SPICE NETLIST
***************************************

.SUBCKT reg1w1 WE RE D CLK Q vss! vdd! Qb
** N=18 EP=8 IP=0 FDC=28
M0 vss! WE 1 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=310 $Y=600 $D=1
M1 4 RE vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=690 $Y=600 $D=1
M2 5 WE D vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=1425 $Y=600 $D=1
M3 vss! 5 12 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=2160 $Y=600 $D=1
M4 6 12 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=1.26e-14 PD=5.25e-07 PS=4.6e-07 $X=2540 $Y=600 $D=1
M5 5 1 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=2985 $Y=600 $D=1
M6 7 RE 6 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.2375e-14 PD=4.55e-07 PS=4.55e-07 $X=3795 $Y=600 $D=1
M7 vss! 9 8 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=4530 $Y=600 $D=1
M8 9 CLK vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=9e-15 AS=1.26e-14 PD=3.8e-07 PS=4.6e-07 $X=4910 $Y=600 $D=1
M9 14 7 vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.5525e-14 AS=9e-15 PD=5.25e-07 PS=3.8e-07 $X=5570 $Y=600 $D=1
M10 10 8 14 vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.2375e-14 AS=1.5525e-14 PD=4.55e-07 PS=5.25e-07 $X=6015 $Y=600 $D=1
M11 vss! 10 Q vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9e-15 PD=4.6e-07 PS=3.8e-07 $X=6750 $Y=600 $D=1
M12 Qb Q vss! vss! NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=7130 $Y=600 $D=1
M13 10 9 Qb vss! NMOS_VTL L=5e-08 W=9e-08 AD=2.4975e-14 AS=1.26e-14 PD=7.35e-07 PS=4.6e-07 $X=7510 $Y=600 $D=1
M14 vdd! WE 1 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=310 $Y=1850 $D=0
M15 4 RE vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=690 $Y=1850 $D=0
M16 5 1 D vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=1425 $Y=1850 $D=0
M17 vdd! 5 12 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=2160 $Y=1850 $D=0
M18 6 12 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=2.52e-14 PD=7.05e-07 PS=6.4e-07 $X=2540 $Y=1850 $D=0
M19 5 WE 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=2985 $Y=1850 $D=0
M20 7 4 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=2.475e-14 PD=6.35e-07 PS=6.35e-07 $X=3795 $Y=1850 $D=0
M21 vdd! 9 8 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=4530 $Y=1850 $D=0
M22 9 CLK vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.8e-14 AS=2.52e-14 PD=5.6e-07 PS=6.4e-07 $X=4910 $Y=1850 $D=0
M23 14 7 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=3.105e-14 AS=1.8e-14 PD=7.05e-07 PS=5.6e-07 $X=5570 $Y=1850 $D=0
M24 10 9 14 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.475e-14 AS=3.105e-14 PD=6.35e-07 PS=7.05e-07 $X=6015 $Y=1850 $D=0
M25 vdd! 10 Q vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.8e-14 PD=6.4e-07 PS=5.6e-07 $X=6750 $Y=1850 $D=0
M26 Qb Q vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=5.58e-14 AS=2.52e-14 PD=9.8e-07 PS=6.4e-07 $X=7130 $Y=1850 $D=0
M27 10 8 Qb vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=5.58e-14 PD=5.75e-07 PS=9.8e-07 $X=7850 $Y=1850 $D=0
.ENDS
***************************************
