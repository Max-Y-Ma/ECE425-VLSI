/home/maxma2/Documents/Coursework/ece425/mp3/lib/stdcells.lef